library verilog;
use verilog.vl_types.all;
entity tb_main is
end tb_main;
