
module myfir ( clk, rst_n, din, vin, b0, b1, b2, b3, b4, b5, b6, b7, b8, b9, 
        b10, dout, vout );
  input [13:0] din;
  input [13:0] b0;
  input [13:0] b1;
  input [13:0] b2;
  input [13:0] b3;
  input [13:0] b4;
  input [13:0] b5;
  input [13:0] b6;
  input [13:0] b7;
  input [13:0] b8;
  input [13:0] b9;
  input [13:0] b10;
  output [13:0] dout;
  input clk, rst_n, vin;
  output vout;
  wire   my_filter_n2, my_filter_q_reg_chain_10__0_,
         my_filter_q_reg_chain_10__1_, my_filter_q_reg_chain_10__2_,
         my_filter_q_reg_chain_10__3_, my_filter_q_reg_chain_10__4_,
         my_filter_q_reg_chain_10__5_, my_filter_q_reg_chain_10__6_,
         my_filter_q_reg_chain_10__7_, my_filter_q_reg_chain_10__8_,
         my_filter_q_reg_chain_10__9_, my_filter_q_reg_chain_10__10_,
         my_filter_q_reg_chain_10__11_, my_filter_q_reg_chain_10__12_,
         my_filter_q_reg_chain_10__13_, my_filter_q_reg_chain_9__0_,
         my_filter_q_reg_chain_9__1_, my_filter_q_reg_chain_9__2_,
         my_filter_q_reg_chain_9__3_, my_filter_q_reg_chain_9__4_,
         my_filter_q_reg_chain_9__5_, my_filter_q_reg_chain_9__6_,
         my_filter_q_reg_chain_9__7_, my_filter_q_reg_chain_9__8_,
         my_filter_q_reg_chain_9__9_, my_filter_q_reg_chain_9__10_,
         my_filter_q_reg_chain_9__11_, my_filter_q_reg_chain_9__12_,
         my_filter_q_reg_chain_9__13_, my_filter_q_reg_chain_8__0_,
         my_filter_q_reg_chain_8__1_, my_filter_q_reg_chain_8__2_,
         my_filter_q_reg_chain_8__3_, my_filter_q_reg_chain_8__4_,
         my_filter_q_reg_chain_8__5_, my_filter_q_reg_chain_8__6_,
         my_filter_q_reg_chain_8__7_, my_filter_q_reg_chain_8__8_,
         my_filter_q_reg_chain_8__9_, my_filter_q_reg_chain_8__10_,
         my_filter_q_reg_chain_8__11_, my_filter_q_reg_chain_8__12_,
         my_filter_q_reg_chain_8__13_, my_filter_q_reg_chain_7__0_,
         my_filter_q_reg_chain_7__1_, my_filter_q_reg_chain_7__2_,
         my_filter_q_reg_chain_7__3_, my_filter_q_reg_chain_7__4_,
         my_filter_q_reg_chain_7__5_, my_filter_q_reg_chain_7__6_,
         my_filter_q_reg_chain_7__7_, my_filter_q_reg_chain_7__8_,
         my_filter_q_reg_chain_7__9_, my_filter_q_reg_chain_7__10_,
         my_filter_q_reg_chain_7__11_, my_filter_q_reg_chain_7__12_,
         my_filter_q_reg_chain_7__13_, my_filter_q_reg_chain_6__0_,
         my_filter_q_reg_chain_6__1_, my_filter_q_reg_chain_6__2_,
         my_filter_q_reg_chain_6__3_, my_filter_q_reg_chain_6__4_,
         my_filter_q_reg_chain_6__5_, my_filter_q_reg_chain_6__6_,
         my_filter_q_reg_chain_6__7_, my_filter_q_reg_chain_6__8_,
         my_filter_q_reg_chain_6__9_, my_filter_q_reg_chain_6__10_,
         my_filter_q_reg_chain_6__11_, my_filter_q_reg_chain_6__12_,
         my_filter_q_reg_chain_6__13_, my_filter_q_reg_chain_5__0_,
         my_filter_q_reg_chain_5__1_, my_filter_q_reg_chain_5__2_,
         my_filter_q_reg_chain_5__3_, my_filter_q_reg_chain_5__4_,
         my_filter_q_reg_chain_5__5_, my_filter_q_reg_chain_5__6_,
         my_filter_q_reg_chain_5__7_, my_filter_q_reg_chain_5__8_,
         my_filter_q_reg_chain_5__9_, my_filter_q_reg_chain_5__10_,
         my_filter_q_reg_chain_5__11_, my_filter_q_reg_chain_5__12_,
         my_filter_q_reg_chain_5__13_, my_filter_q_reg_chain_4__0_,
         my_filter_q_reg_chain_4__1_, my_filter_q_reg_chain_4__2_,
         my_filter_q_reg_chain_4__3_, my_filter_q_reg_chain_4__4_,
         my_filter_q_reg_chain_4__5_, my_filter_q_reg_chain_4__6_,
         my_filter_q_reg_chain_4__7_, my_filter_q_reg_chain_4__8_,
         my_filter_q_reg_chain_4__9_, my_filter_q_reg_chain_4__10_,
         my_filter_q_reg_chain_4__11_, my_filter_q_reg_chain_4__12_,
         my_filter_q_reg_chain_4__13_, my_filter_q_reg_chain_3__0_,
         my_filter_q_reg_chain_3__1_, my_filter_q_reg_chain_3__2_,
         my_filter_q_reg_chain_3__3_, my_filter_q_reg_chain_3__4_,
         my_filter_q_reg_chain_3__5_, my_filter_q_reg_chain_3__6_,
         my_filter_q_reg_chain_3__7_, my_filter_q_reg_chain_3__8_,
         my_filter_q_reg_chain_3__9_, my_filter_q_reg_chain_3__10_,
         my_filter_q_reg_chain_3__11_, my_filter_q_reg_chain_3__12_,
         my_filter_q_reg_chain_3__13_, my_filter_q_reg_chain_2__0_,
         my_filter_q_reg_chain_2__1_, my_filter_q_reg_chain_2__2_,
         my_filter_q_reg_chain_2__3_, my_filter_q_reg_chain_2__4_,
         my_filter_q_reg_chain_2__5_, my_filter_q_reg_chain_2__6_,
         my_filter_q_reg_chain_2__7_, my_filter_q_reg_chain_2__8_,
         my_filter_q_reg_chain_2__9_, my_filter_q_reg_chain_2__10_,
         my_filter_q_reg_chain_2__11_, my_filter_q_reg_chain_2__12_,
         my_filter_q_reg_chain_2__13_, my_filter_q_reg_chain_1__0_,
         my_filter_q_reg_chain_1__1_, my_filter_q_reg_chain_1__2_,
         my_filter_q_reg_chain_1__3_, my_filter_q_reg_chain_1__4_,
         my_filter_q_reg_chain_1__5_, my_filter_q_reg_chain_1__6_,
         my_filter_q_reg_chain_1__7_, my_filter_q_reg_chain_1__8_,
         my_filter_q_reg_chain_1__9_, my_filter_q_reg_chain_1__10_,
         my_filter_q_reg_chain_1__11_, my_filter_q_reg_chain_1__12_,
         my_filter_q_reg_chain_1__13_, my_filter_en_reg_out,
         my_filter_q_reg_samp_0_, my_filter_q_reg_samp_1_,
         my_filter_q_reg_samp_2_, my_filter_q_reg_samp_3_,
         my_filter_q_reg_samp_4_, my_filter_q_reg_samp_5_,
         my_filter_q_reg_samp_6_, my_filter_q_reg_samp_7_,
         my_filter_q_reg_samp_8_, my_filter_q_reg_samp_9_,
         my_filter_q_reg_samp_10_, my_filter_q_reg_samp_11_,
         my_filter_q_reg_samp_12_, my_filter_q_reg_samp_13_,
         my_filter_reg_samples_n46, my_filter_reg_samples_n45,
         my_filter_reg_samples_n44, my_filter_reg_samples_n43,
         my_filter_reg_samples_n42, my_filter_reg_samples_n41,
         my_filter_reg_samples_n40, my_filter_reg_samples_n39,
         my_filter_reg_samples_n38, my_filter_reg_samples_n37,
         my_filter_reg_samples_n36, my_filter_reg_samples_n35,
         my_filter_reg_samples_n34, my_filter_reg_samples_n33,
         my_filter_reg_samples_n32, my_filter_reg_samples_n31,
         my_filter_reg_samples_n30, my_filter_reg_samples_n29,
         my_filter_reg_samples_n28, my_filter_reg_samples_n27,
         my_filter_reg_samples_n26, my_filter_reg_samples_n25,
         my_filter_reg_samples_n24, my_filter_reg_samples_n23,
         my_filter_reg_samples_n22, my_filter_reg_samples_n21,
         my_filter_reg_samples_n20, my_filter_reg_samples_n19,
         my_filter_reg_samples_n18, my_filter_reg_samples_n17,
         my_filter_reg_samples_n16, my_filter_reg_samples_n15,
         my_filter_reg_samples_n14, my_filter_reg_samples_n13,
         my_filter_reg_samples_n12, my_filter_reg_samples_n11,
         my_filter_reg_samples_n10, my_filter_reg_samples_n9,
         my_filter_reg_samples_n8, my_filter_reg_samples_n7,
         my_filter_reg_samples_n6, my_filter_reg_samples_n5,
         my_filter_reg_samples_n4, my_filter_reg_samples_n3,
         my_filter_reg_samples_n2, my_filter_reg_coefficients_n505,
         my_filter_reg_coefficients_n504, my_filter_reg_coefficients_n503,
         my_filter_reg_coefficients_n502, my_filter_reg_coefficients_n501,
         my_filter_reg_coefficients_n500, my_filter_reg_coefficients_n499,
         my_filter_reg_coefficients_n498, my_filter_reg_coefficients_n497,
         my_filter_reg_coefficients_n496, my_filter_reg_coefficients_n495,
         my_filter_reg_coefficients_n494, my_filter_reg_coefficients_n493,
         my_filter_reg_coefficients_n492, my_filter_reg_coefficients_n491,
         my_filter_reg_coefficients_n490, my_filter_reg_coefficients_n489,
         my_filter_reg_coefficients_n488, my_filter_reg_coefficients_n487,
         my_filter_reg_coefficients_n486, my_filter_reg_coefficients_n485,
         my_filter_reg_coefficients_n484, my_filter_reg_coefficients_n483,
         my_filter_reg_coefficients_n482, my_filter_reg_coefficients_n481,
         my_filter_reg_coefficients_n480, my_filter_reg_coefficients_n479,
         my_filter_reg_coefficients_n478, my_filter_reg_coefficients_n477,
         my_filter_reg_coefficients_n476, my_filter_reg_coefficients_n475,
         my_filter_reg_coefficients_n474, my_filter_reg_coefficients_n473,
         my_filter_reg_coefficients_n472, my_filter_reg_coefficients_n471,
         my_filter_reg_coefficients_n470, my_filter_reg_coefficients_n469,
         my_filter_reg_coefficients_n468, my_filter_reg_coefficients_n467,
         my_filter_reg_coefficients_n466, my_filter_reg_coefficients_n465,
         my_filter_reg_coefficients_n464, my_filter_reg_coefficients_n463,
         my_filter_reg_coefficients_n462, my_filter_reg_coefficients_n461,
         my_filter_reg_coefficients_n460, my_filter_reg_coefficients_n459,
         my_filter_reg_coefficients_n458, my_filter_reg_coefficients_n457,
         my_filter_reg_coefficients_n456, my_filter_reg_coefficients_n455,
         my_filter_reg_coefficients_n454, my_filter_reg_coefficients_n453,
         my_filter_reg_coefficients_n452, my_filter_reg_coefficients_n451,
         my_filter_reg_coefficients_n450, my_filter_reg_coefficients_n449,
         my_filter_reg_coefficients_n448, my_filter_reg_coefficients_n447,
         my_filter_reg_coefficients_n446, my_filter_reg_coefficients_n445,
         my_filter_reg_coefficients_n444, my_filter_reg_coefficients_n443,
         my_filter_reg_coefficients_n442, my_filter_reg_coefficients_n441,
         my_filter_reg_coefficients_n440, my_filter_reg_coefficients_n439,
         my_filter_reg_coefficients_n438, my_filter_reg_coefficients_n437,
         my_filter_reg_coefficients_n436, my_filter_reg_coefficients_n435,
         my_filter_reg_coefficients_n434, my_filter_reg_coefficients_n433,
         my_filter_reg_coefficients_n432, my_filter_reg_coefficients_n431,
         my_filter_reg_coefficients_n430, my_filter_reg_coefficients_n429,
         my_filter_reg_coefficients_n428, my_filter_reg_coefficients_n427,
         my_filter_reg_coefficients_n426, my_filter_reg_coefficients_n425,
         my_filter_reg_coefficients_n424, my_filter_reg_coefficients_n423,
         my_filter_reg_coefficients_n422, my_filter_reg_coefficients_n421,
         my_filter_reg_coefficients_n420, my_filter_reg_coefficients_n419,
         my_filter_reg_coefficients_n418, my_filter_reg_coefficients_n417,
         my_filter_reg_coefficients_n416, my_filter_reg_coefficients_n415,
         my_filter_reg_coefficients_n414, my_filter_reg_coefficients_n413,
         my_filter_reg_coefficients_n412, my_filter_reg_coefficients_n411,
         my_filter_reg_coefficients_n410, my_filter_reg_coefficients_n409,
         my_filter_reg_coefficients_n408, my_filter_reg_coefficients_n407,
         my_filter_reg_coefficients_n406, my_filter_reg_coefficients_n405,
         my_filter_reg_coefficients_n404, my_filter_reg_coefficients_n403,
         my_filter_reg_coefficients_n402, my_filter_reg_coefficients_n401,
         my_filter_reg_coefficients_n400, my_filter_reg_coefficients_n399,
         my_filter_reg_coefficients_n398, my_filter_reg_coefficients_n397,
         my_filter_reg_coefficients_n396, my_filter_reg_coefficients_n395,
         my_filter_reg_coefficients_n394, my_filter_reg_coefficients_n393,
         my_filter_reg_coefficients_n392, my_filter_reg_coefficients_n391,
         my_filter_reg_coefficients_n390, my_filter_reg_coefficients_n389,
         my_filter_reg_coefficients_n388, my_filter_reg_coefficients_n387,
         my_filter_reg_coefficients_n386, my_filter_reg_coefficients_n385,
         my_filter_reg_coefficients_n384, my_filter_reg_coefficients_n383,
         my_filter_reg_coefficients_n382, my_filter_reg_coefficients_n381,
         my_filter_reg_coefficients_n380, my_filter_reg_coefficients_n379,
         my_filter_reg_coefficients_n378, my_filter_reg_coefficients_n377,
         my_filter_reg_coefficients_n376, my_filter_reg_coefficients_n375,
         my_filter_reg_coefficients_n374, my_filter_reg_coefficients_n373,
         my_filter_reg_coefficients_n372, my_filter_reg_coefficients_n371,
         my_filter_reg_coefficients_n370, my_filter_reg_coefficients_n369,
         my_filter_reg_coefficients_n368, my_filter_reg_coefficients_n367,
         my_filter_reg_coefficients_n366, my_filter_reg_coefficients_n365,
         my_filter_reg_coefficients_n364, my_filter_reg_coefficients_n363,
         my_filter_reg_coefficients_n362, my_filter_reg_coefficients_n361,
         my_filter_reg_coefficients_n360, my_filter_reg_coefficients_n359,
         my_filter_reg_coefficients_n358, my_filter_reg_coefficients_n357,
         my_filter_reg_coefficients_n356, my_filter_reg_coefficients_n355,
         my_filter_reg_coefficients_n354, my_filter_reg_coefficients_n353,
         my_filter_reg_coefficients_n352, my_filter_reg_coefficients_n351,
         my_filter_reg_coefficients_n350, my_filter_reg_coefficients_n349,
         my_filter_reg_coefficients_n348, my_filter_reg_coefficients_n347,
         my_filter_reg_coefficients_n346, my_filter_reg_coefficients_n345,
         my_filter_reg_coefficients_n344, my_filter_reg_coefficients_n343,
         my_filter_reg_coefficients_n342, my_filter_reg_coefficients_n341,
         my_filter_reg_coefficients_n340, my_filter_reg_coefficients_n339,
         my_filter_reg_coefficients_n338, my_filter_reg_coefficients_n337,
         my_filter_reg_coefficients_n336, my_filter_reg_coefficients_n335,
         my_filter_reg_coefficients_n334, my_filter_reg_coefficients_n333,
         my_filter_reg_coefficients_n332, my_filter_reg_coefficients_n331,
         my_filter_reg_coefficients_n330, my_filter_reg_coefficients_n329,
         my_filter_reg_coefficients_n328, my_filter_reg_coefficients_n327,
         my_filter_reg_coefficients_n326, my_filter_reg_coefficients_n325,
         my_filter_reg_coefficients_n324, my_filter_reg_coefficients_n323,
         my_filter_reg_coefficients_n322, my_filter_reg_coefficients_n321,
         my_filter_reg_coefficients_n320, my_filter_reg_coefficients_n319,
         my_filter_reg_coefficients_n318, my_filter_reg_coefficients_n317,
         my_filter_reg_coefficients_n316, my_filter_reg_coefficients_n315,
         my_filter_reg_coefficients_n314, my_filter_reg_coefficients_n313,
         my_filter_reg_coefficients_n312, my_filter_reg_coefficients_n311,
         my_filter_reg_coefficients_n310, my_filter_reg_coefficients_n309,
         my_filter_reg_coefficients_n308, my_filter_reg_coefficients_n307,
         my_filter_reg_coefficients_n306, my_filter_reg_coefficients_n305,
         my_filter_reg_coefficients_n304, my_filter_reg_coefficients_n303,
         my_filter_reg_coefficients_n302, my_filter_reg_coefficients_n301,
         my_filter_reg_coefficients_n300, my_filter_reg_coefficients_n299,
         my_filter_reg_coefficients_n298, my_filter_reg_coefficients_n297,
         my_filter_reg_coefficients_n296, my_filter_reg_coefficients_n295,
         my_filter_reg_coefficients_n294, my_filter_reg_coefficients_n293,
         my_filter_reg_coefficients_n292, my_filter_reg_coefficients_n291,
         my_filter_reg_coefficients_n290, my_filter_reg_coefficients_n289,
         my_filter_reg_coefficients_n288, my_filter_reg_coefficients_n287,
         my_filter_reg_coefficients_n286, my_filter_reg_coefficients_n285,
         my_filter_reg_coefficients_n284, my_filter_reg_coefficients_n283,
         my_filter_reg_coefficients_n282, my_filter_reg_coefficients_n281,
         my_filter_reg_coefficients_n280, my_filter_reg_coefficients_n279,
         my_filter_reg_coefficients_n278, my_filter_reg_coefficients_n277,
         my_filter_reg_coefficients_n276, my_filter_reg_coefficients_n275,
         my_filter_reg_coefficients_n274, my_filter_reg_coefficients_n273,
         my_filter_reg_coefficients_n272, my_filter_reg_coefficients_n271,
         my_filter_reg_coefficients_n270, my_filter_reg_coefficients_n269,
         my_filter_reg_coefficients_n268, my_filter_reg_coefficients_n267,
         my_filter_reg_coefficients_n266, my_filter_reg_coefficients_n265,
         my_filter_reg_coefficients_n264, my_filter_reg_coefficients_n263,
         my_filter_reg_coefficients_n262, my_filter_reg_coefficients_n261,
         my_filter_reg_coefficients_n260, my_filter_reg_coefficients_n259,
         my_filter_reg_coefficients_n258, my_filter_reg_coefficients_n257,
         my_filter_reg_coefficients_n256, my_filter_reg_coefficients_n255,
         my_filter_reg_coefficients_n254, my_filter_reg_coefficients_n253,
         my_filter_reg_coefficients_n252, my_filter_reg_coefficients_n251,
         my_filter_reg_coefficients_n250, my_filter_reg_coefficients_n249,
         my_filter_reg_coefficients_n248, my_filter_reg_coefficients_n247,
         my_filter_reg_coefficients_n246, my_filter_reg_coefficients_n245,
         my_filter_reg_coefficients_n244, my_filter_reg_coefficients_n243,
         my_filter_reg_coefficients_n242, my_filter_reg_coefficients_n241,
         my_filter_reg_coefficients_n240, my_filter_reg_coefficients_n239,
         my_filter_reg_coefficients_n238, my_filter_reg_coefficients_n237,
         my_filter_reg_coefficients_n236, my_filter_reg_coefficients_n235,
         my_filter_reg_coefficients_n234, my_filter_reg_coefficients_n233,
         my_filter_reg_coefficients_n232, my_filter_reg_coefficients_n231,
         my_filter_reg_coefficients_n230, my_filter_reg_coefficients_n229,
         my_filter_reg_coefficients_n228, my_filter_reg_coefficients_n227,
         my_filter_reg_coefficients_n226, my_filter_reg_coefficients_n225,
         my_filter_reg_coefficients_n224, my_filter_reg_coefficients_n223,
         my_filter_reg_coefficients_n222, my_filter_reg_coefficients_n221,
         my_filter_reg_coefficients_n220, my_filter_reg_coefficients_n219,
         my_filter_reg_coefficients_n218, my_filter_reg_coefficients_n217,
         my_filter_reg_coefficients_n216, my_filter_reg_coefficients_n215,
         my_filter_reg_coefficients_n214, my_filter_reg_coefficients_n213,
         my_filter_reg_coefficients_n212, my_filter_reg_coefficients_n211,
         my_filter_reg_coefficients_n210, my_filter_reg_coefficients_n209,
         my_filter_reg_coefficients_n208, my_filter_reg_coefficients_n207,
         my_filter_reg_coefficients_n206, my_filter_reg_coefficients_n205,
         my_filter_reg_coefficients_n204, my_filter_reg_coefficients_n203,
         my_filter_reg_coefficients_n202, my_filter_reg_coefficients_n201,
         my_filter_reg_coefficients_n200, my_filter_reg_coefficients_n199,
         my_filter_reg_coefficients_n198, my_filter_reg_coefficients_n197,
         my_filter_reg_coefficients_n196, my_filter_reg_coefficients_n195,
         my_filter_reg_coefficients_n194, my_filter_reg_coefficients_n193,
         my_filter_reg_coefficients_n192, my_filter_reg_coefficients_n191,
         my_filter_reg_coefficients_n190, my_filter_reg_coefficients_n189,
         my_filter_reg_coefficients_n188, my_filter_reg_coefficients_n187,
         my_filter_reg_coefficients_n186, my_filter_reg_coefficients_n185,
         my_filter_reg_coefficients_n184, my_filter_reg_coefficients_n183,
         my_filter_reg_coefficients_n182, my_filter_reg_coefficients_n181,
         my_filter_reg_coefficients_n180, my_filter_reg_coefficients_n179,
         my_filter_reg_coefficients_n178, my_filter_reg_coefficients_n177,
         my_filter_reg_coefficients_n176, my_filter_reg_coefficients_n175,
         my_filter_reg_coefficients_n174, my_filter_reg_coefficients_n173,
         my_filter_reg_coefficients_n172, my_filter_reg_coefficients_n171,
         my_filter_reg_coefficients_n170, my_filter_reg_coefficients_n169,
         my_filter_reg_coefficients_n168, my_filter_reg_coefficients_n167,
         my_filter_reg_coefficients_n166, my_filter_reg_coefficients_n165,
         my_filter_reg_coefficients_n164, my_filter_reg_coefficients_n163,
         my_filter_reg_coefficients_n162, my_filter_reg_coefficients_n161,
         my_filter_reg_coefficients_n160, my_filter_reg_coefficients_n159,
         my_filter_reg_coefficients_n158, my_filter_reg_coefficients_n157,
         my_filter_reg_coefficients_n156, my_filter_reg_coefficients_n155,
         my_filter_reg_coefficients_n154, my_filter_reg_coefficients_n153,
         my_filter_reg_coefficients_n152, my_filter_reg_coefficients_n151,
         my_filter_reg_coefficients_n150, my_filter_reg_coefficients_n149,
         my_filter_reg_coefficients_n148, my_filter_reg_coefficients_n147,
         my_filter_reg_coefficients_n146, my_filter_reg_coefficients_n145,
         my_filter_reg_coefficients_n144, my_filter_reg_coefficients_n143,
         my_filter_reg_coefficients_n142, my_filter_reg_coefficients_n141,
         my_filter_reg_coefficients_n140, my_filter_reg_coefficients_n139,
         my_filter_reg_coefficients_n138, my_filter_reg_coefficients_n137,
         my_filter_reg_coefficients_n136, my_filter_reg_coefficients_n135,
         my_filter_reg_coefficients_n134, my_filter_reg_coefficients_n133,
         my_filter_reg_coefficients_n132, my_filter_reg_coefficients_n131,
         my_filter_reg_coefficients_n130, my_filter_reg_coefficients_n129,
         my_filter_reg_coefficients_n128, my_filter_reg_coefficients_n127,
         my_filter_reg_coefficients_n126, my_filter_reg_coefficients_n125,
         my_filter_reg_coefficients_n124, my_filter_reg_coefficients_n123,
         my_filter_reg_coefficients_n122, my_filter_reg_coefficients_n121,
         my_filter_reg_coefficients_n120, my_filter_reg_coefficients_n119,
         my_filter_reg_coefficients_n118, my_filter_reg_coefficients_n117,
         my_filter_reg_coefficients_n116, my_filter_reg_coefficients_n115,
         my_filter_reg_coefficients_n114, my_filter_reg_coefficients_n113,
         my_filter_reg_coefficients_n112, my_filter_reg_coefficients_n111,
         my_filter_reg_coefficients_n110, my_filter_reg_coefficients_n109,
         my_filter_reg_coefficients_n108, my_filter_reg_coefficients_n107,
         my_filter_reg_coefficients_n106, my_filter_reg_coefficients_n105,
         my_filter_reg_coefficients_n104, my_filter_reg_coefficients_n103,
         my_filter_reg_coefficients_n102, my_filter_reg_coefficients_n101,
         my_filter_reg_coefficients_n100, my_filter_reg_coefficients_n99,
         my_filter_reg_coefficients_n98, my_filter_reg_coefficients_n97,
         my_filter_reg_coefficients_n96, my_filter_reg_coefficients_n95,
         my_filter_reg_coefficients_n94, my_filter_reg_coefficients_n93,
         my_filter_reg_coefficients_n92, my_filter_reg_coefficients_n91,
         my_filter_reg_coefficients_n90, my_filter_reg_coefficients_n89,
         my_filter_reg_coefficients_n88, my_filter_reg_coefficients_n87,
         my_filter_reg_coefficients_n86, my_filter_reg_coefficients_n85,
         my_filter_reg_coefficients_n84, my_filter_reg_coefficients_n83,
         my_filter_reg_coefficients_n82, my_filter_reg_coefficients_n81,
         my_filter_reg_coefficients_n80, my_filter_reg_coefficients_n79,
         my_filter_reg_coefficients_n78, my_filter_reg_coefficients_n77,
         my_filter_reg_coefficients_n76, my_filter_reg_coefficients_n75,
         my_filter_reg_coefficients_n74, my_filter_reg_coefficients_n73,
         my_filter_reg_coefficients_n72, my_filter_reg_coefficients_n71,
         my_filter_reg_coefficients_n70, my_filter_reg_coefficients_n69,
         my_filter_reg_coefficients_n68, my_filter_reg_coefficients_n67,
         my_filter_reg_coefficients_n66, my_filter_reg_coefficients_n65,
         my_filter_reg_coefficients_n64, my_filter_reg_coefficients_n63,
         my_filter_reg_coefficients_n62, my_filter_reg_coefficients_n61,
         my_filter_reg_coefficients_n60, my_filter_reg_coefficients_n59,
         my_filter_reg_coefficients_n58, my_filter_reg_coefficients_n57,
         my_filter_reg_coefficients_n56, my_filter_reg_coefficients_n55,
         my_filter_reg_coefficients_n54, my_filter_reg_coefficients_n53,
         my_filter_reg_coefficients_n52, my_filter_reg_coefficients_n51,
         my_filter_reg_coefficients_n50, my_filter_reg_coefficients_n49,
         my_filter_reg_coefficients_n48, my_filter_reg_coefficients_n47,
         my_filter_reg_coefficients_n46, my_filter_reg_coefficients_n45,
         my_filter_reg_coefficients_n44, my_filter_reg_coefficients_n43,
         my_filter_reg_coefficients_n42, my_filter_reg_coefficients_n41,
         my_filter_reg_coefficients_n40, my_filter_reg_coefficients_n39,
         my_filter_reg_coefficients_n38, my_filter_reg_coefficients_n37,
         my_filter_reg_coefficients_n36, my_filter_reg_coefficients_n35,
         my_filter_reg_coefficients_n34, my_filter_reg_coefficients_n33,
         my_filter_reg_coefficients_n32, my_filter_reg_coefficients_n31,
         my_filter_reg_coefficients_n30, my_filter_reg_coefficients_n29,
         my_filter_reg_coefficients_n28, my_filter_reg_coefficients_n27,
         my_filter_reg_coefficients_n26, my_filter_reg_coefficients_n25,
         my_filter_reg_coefficients_n24, my_filter_reg_coefficients_n23,
         my_filter_reg_coefficients_n22, my_filter_reg_coefficients_n21,
         my_filter_reg_coefficients_n20, my_filter_reg_coefficients_n19,
         my_filter_reg_coefficients_n18, my_filter_reg_coefficients_n17,
         my_filter_reg_coefficients_n16, my_filter_reg_coefficients_n15,
         my_filter_reg_coefficients_n14, my_filter_reg_coefficients_n13,
         my_filter_reg_coefficients_n12, my_filter_reg_coefficients_n11,
         my_filter_reg_coefficients_n10, my_filter_reg_coefficients_n9,
         my_filter_reg_coefficients_n8, my_filter_reg_coefficients_n7,
         my_filter_reg_coefficients_n6, my_filter_reg_coefficients_n5,
         my_filter_reg_coefficients_n4, my_filter_reg_coefficients_n3,
         my_filter_reg_coefficients_n2, my_filter_reg_out_n47,
         my_filter_reg_out_n46, my_filter_reg_out_n44, my_filter_reg_out_n43,
         my_filter_reg_out_n42, my_filter_reg_out_n41, my_filter_reg_out_n40,
         my_filter_reg_out_n39, my_filter_reg_out_n38, my_filter_reg_out_n37,
         my_filter_reg_out_n36, my_filter_reg_out_n35, my_filter_reg_out_n34,
         my_filter_reg_out_n33, my_filter_reg_out_n32, my_filter_reg_out_n31,
         my_filter_reg_out_n30, my_filter_reg_out_n29, my_filter_reg_out_n28,
         my_filter_reg_out_n27, my_filter_reg_out_n26, my_filter_reg_out_n25,
         my_filter_reg_out_n24, my_filter_reg_out_n23, my_filter_reg_out_n22,
         my_filter_reg_out_n21, my_filter_reg_out_n20, my_filter_reg_out_n19,
         my_filter_reg_out_n18, my_filter_reg_out_n17, my_filter_reg_out_n16,
         my_filter_reg_out_n15, my_filter_reg_out_n14, my_filter_reg_out_n13,
         my_filter_reg_out_n12, my_filter_reg_out_n11, my_filter_reg_out_n10,
         my_filter_reg_out_n9, my_filter_reg_out_n8, my_filter_reg_out_n7,
         my_filter_reg_out_n6, my_filter_reg_out_n5, my_filter_reg_out_n4,
         my_filter_reg_out_n3, my_filter_reg_out_n2, my_filter_delay_line_n15,
         my_filter_delay_line_n14, my_filter_delay_line_n13,
         my_filter_delay_line_n12, my_filter_delay_line_n11,
         my_filter_delay_line_n10, my_filter_delay_line_n9,
         my_filter_delay_line_n8, my_filter_delay_line_delay_chain_0_n50,
         my_filter_delay_line_delay_chain_0_n49,
         my_filter_delay_line_delay_chain_0_n48,
         my_filter_delay_line_delay_chain_0_n44,
         my_filter_delay_line_delay_chain_0_n43,
         my_filter_delay_line_delay_chain_0_n42,
         my_filter_delay_line_delay_chain_0_n41,
         my_filter_delay_line_delay_chain_0_n40,
         my_filter_delay_line_delay_chain_0_n39,
         my_filter_delay_line_delay_chain_0_n38,
         my_filter_delay_line_delay_chain_0_n37,
         my_filter_delay_line_delay_chain_0_n36,
         my_filter_delay_line_delay_chain_0_n35,
         my_filter_delay_line_delay_chain_0_n34,
         my_filter_delay_line_delay_chain_0_n33,
         my_filter_delay_line_delay_chain_0_n32,
         my_filter_delay_line_delay_chain_0_n31,
         my_filter_delay_line_delay_chain_0_n30,
         my_filter_delay_line_delay_chain_0_n29,
         my_filter_delay_line_delay_chain_0_n28,
         my_filter_delay_line_delay_chain_0_n27,
         my_filter_delay_line_delay_chain_0_n26,
         my_filter_delay_line_delay_chain_0_n25,
         my_filter_delay_line_delay_chain_0_n24,
         my_filter_delay_line_delay_chain_0_n23,
         my_filter_delay_line_delay_chain_0_n22,
         my_filter_delay_line_delay_chain_0_n21,
         my_filter_delay_line_delay_chain_0_n20,
         my_filter_delay_line_delay_chain_0_n19,
         my_filter_delay_line_delay_chain_0_n18,
         my_filter_delay_line_delay_chain_0_n17,
         my_filter_delay_line_delay_chain_0_n16,
         my_filter_delay_line_delay_chain_0_n15,
         my_filter_delay_line_delay_chain_0_n14,
         my_filter_delay_line_delay_chain_0_n13,
         my_filter_delay_line_delay_chain_0_n12,
         my_filter_delay_line_delay_chain_0_n11,
         my_filter_delay_line_delay_chain_0_n10,
         my_filter_delay_line_delay_chain_0_n9,
         my_filter_delay_line_delay_chain_0_n8,
         my_filter_delay_line_delay_chain_0_n7,
         my_filter_delay_line_delay_chain_0_n6,
         my_filter_delay_line_delay_chain_0_n5,
         my_filter_delay_line_delay_chain_0_n4,
         my_filter_delay_line_delay_chain_0_n3,
         my_filter_delay_line_delay_chain_0_n2,
         my_filter_delay_line_delay_chain_1_n94,
         my_filter_delay_line_delay_chain_1_n93,
         my_filter_delay_line_delay_chain_1_n92,
         my_filter_delay_line_delay_chain_1_n91,
         my_filter_delay_line_delay_chain_1_n90,
         my_filter_delay_line_delay_chain_1_n89,
         my_filter_delay_line_delay_chain_1_n88,
         my_filter_delay_line_delay_chain_1_n87,
         my_filter_delay_line_delay_chain_1_n86,
         my_filter_delay_line_delay_chain_1_n85,
         my_filter_delay_line_delay_chain_1_n84,
         my_filter_delay_line_delay_chain_1_n83,
         my_filter_delay_line_delay_chain_1_n82,
         my_filter_delay_line_delay_chain_1_n81,
         my_filter_delay_line_delay_chain_1_n80,
         my_filter_delay_line_delay_chain_1_n79,
         my_filter_delay_line_delay_chain_1_n78,
         my_filter_delay_line_delay_chain_1_n77,
         my_filter_delay_line_delay_chain_1_n76,
         my_filter_delay_line_delay_chain_1_n75,
         my_filter_delay_line_delay_chain_1_n74,
         my_filter_delay_line_delay_chain_1_n73,
         my_filter_delay_line_delay_chain_1_n72,
         my_filter_delay_line_delay_chain_1_n71,
         my_filter_delay_line_delay_chain_1_n70,
         my_filter_delay_line_delay_chain_1_n69,
         my_filter_delay_line_delay_chain_1_n68,
         my_filter_delay_line_delay_chain_1_n67,
         my_filter_delay_line_delay_chain_1_n66,
         my_filter_delay_line_delay_chain_1_n65,
         my_filter_delay_line_delay_chain_1_n64,
         my_filter_delay_line_delay_chain_1_n63,
         my_filter_delay_line_delay_chain_1_n62,
         my_filter_delay_line_delay_chain_1_n61,
         my_filter_delay_line_delay_chain_1_n60,
         my_filter_delay_line_delay_chain_1_n59,
         my_filter_delay_line_delay_chain_1_n58,
         my_filter_delay_line_delay_chain_1_n57,
         my_filter_delay_line_delay_chain_1_n56,
         my_filter_delay_line_delay_chain_1_n55,
         my_filter_delay_line_delay_chain_1_n54,
         my_filter_delay_line_delay_chain_1_n53,
         my_filter_delay_line_delay_chain_1_n52,
         my_filter_delay_line_delay_chain_1_n51,
         my_filter_delay_line_delay_chain_1_n50,
         my_filter_delay_line_delay_chain_1_n49,
         my_filter_delay_line_delay_chain_1_n48,
         my_filter_delay_line_delay_chain_2_n94,
         my_filter_delay_line_delay_chain_2_n93,
         my_filter_delay_line_delay_chain_2_n92,
         my_filter_delay_line_delay_chain_2_n91,
         my_filter_delay_line_delay_chain_2_n90,
         my_filter_delay_line_delay_chain_2_n89,
         my_filter_delay_line_delay_chain_2_n88,
         my_filter_delay_line_delay_chain_2_n87,
         my_filter_delay_line_delay_chain_2_n86,
         my_filter_delay_line_delay_chain_2_n85,
         my_filter_delay_line_delay_chain_2_n84,
         my_filter_delay_line_delay_chain_2_n83,
         my_filter_delay_line_delay_chain_2_n82,
         my_filter_delay_line_delay_chain_2_n81,
         my_filter_delay_line_delay_chain_2_n80,
         my_filter_delay_line_delay_chain_2_n79,
         my_filter_delay_line_delay_chain_2_n78,
         my_filter_delay_line_delay_chain_2_n77,
         my_filter_delay_line_delay_chain_2_n76,
         my_filter_delay_line_delay_chain_2_n75,
         my_filter_delay_line_delay_chain_2_n74,
         my_filter_delay_line_delay_chain_2_n73,
         my_filter_delay_line_delay_chain_2_n72,
         my_filter_delay_line_delay_chain_2_n71,
         my_filter_delay_line_delay_chain_2_n70,
         my_filter_delay_line_delay_chain_2_n69,
         my_filter_delay_line_delay_chain_2_n68,
         my_filter_delay_line_delay_chain_2_n67,
         my_filter_delay_line_delay_chain_2_n66,
         my_filter_delay_line_delay_chain_2_n65,
         my_filter_delay_line_delay_chain_2_n64,
         my_filter_delay_line_delay_chain_2_n63,
         my_filter_delay_line_delay_chain_2_n62,
         my_filter_delay_line_delay_chain_2_n61,
         my_filter_delay_line_delay_chain_2_n60,
         my_filter_delay_line_delay_chain_2_n59,
         my_filter_delay_line_delay_chain_2_n58,
         my_filter_delay_line_delay_chain_2_n57,
         my_filter_delay_line_delay_chain_2_n56,
         my_filter_delay_line_delay_chain_2_n55,
         my_filter_delay_line_delay_chain_2_n54,
         my_filter_delay_line_delay_chain_2_n53,
         my_filter_delay_line_delay_chain_2_n52,
         my_filter_delay_line_delay_chain_2_n51,
         my_filter_delay_line_delay_chain_2_n50,
         my_filter_delay_line_delay_chain_2_n49,
         my_filter_delay_line_delay_chain_2_n48,
         my_filter_delay_line_delay_chain_3_n94,
         my_filter_delay_line_delay_chain_3_n93,
         my_filter_delay_line_delay_chain_3_n92,
         my_filter_delay_line_delay_chain_3_n91,
         my_filter_delay_line_delay_chain_3_n90,
         my_filter_delay_line_delay_chain_3_n89,
         my_filter_delay_line_delay_chain_3_n88,
         my_filter_delay_line_delay_chain_3_n87,
         my_filter_delay_line_delay_chain_3_n86,
         my_filter_delay_line_delay_chain_3_n85,
         my_filter_delay_line_delay_chain_3_n84,
         my_filter_delay_line_delay_chain_3_n83,
         my_filter_delay_line_delay_chain_3_n82,
         my_filter_delay_line_delay_chain_3_n81,
         my_filter_delay_line_delay_chain_3_n80,
         my_filter_delay_line_delay_chain_3_n79,
         my_filter_delay_line_delay_chain_3_n78,
         my_filter_delay_line_delay_chain_3_n77,
         my_filter_delay_line_delay_chain_3_n76,
         my_filter_delay_line_delay_chain_3_n75,
         my_filter_delay_line_delay_chain_3_n74,
         my_filter_delay_line_delay_chain_3_n73,
         my_filter_delay_line_delay_chain_3_n72,
         my_filter_delay_line_delay_chain_3_n71,
         my_filter_delay_line_delay_chain_3_n70,
         my_filter_delay_line_delay_chain_3_n69,
         my_filter_delay_line_delay_chain_3_n68,
         my_filter_delay_line_delay_chain_3_n67,
         my_filter_delay_line_delay_chain_3_n66,
         my_filter_delay_line_delay_chain_3_n65,
         my_filter_delay_line_delay_chain_3_n64,
         my_filter_delay_line_delay_chain_3_n63,
         my_filter_delay_line_delay_chain_3_n62,
         my_filter_delay_line_delay_chain_3_n61,
         my_filter_delay_line_delay_chain_3_n60,
         my_filter_delay_line_delay_chain_3_n59,
         my_filter_delay_line_delay_chain_3_n58,
         my_filter_delay_line_delay_chain_3_n57,
         my_filter_delay_line_delay_chain_3_n56,
         my_filter_delay_line_delay_chain_3_n55,
         my_filter_delay_line_delay_chain_3_n54,
         my_filter_delay_line_delay_chain_3_n53,
         my_filter_delay_line_delay_chain_3_n52,
         my_filter_delay_line_delay_chain_3_n51,
         my_filter_delay_line_delay_chain_3_n50,
         my_filter_delay_line_delay_chain_3_n49,
         my_filter_delay_line_delay_chain_3_n48,
         my_filter_delay_line_delay_chain_4_n94,
         my_filter_delay_line_delay_chain_4_n93,
         my_filter_delay_line_delay_chain_4_n92,
         my_filter_delay_line_delay_chain_4_n91,
         my_filter_delay_line_delay_chain_4_n90,
         my_filter_delay_line_delay_chain_4_n89,
         my_filter_delay_line_delay_chain_4_n88,
         my_filter_delay_line_delay_chain_4_n87,
         my_filter_delay_line_delay_chain_4_n86,
         my_filter_delay_line_delay_chain_4_n85,
         my_filter_delay_line_delay_chain_4_n84,
         my_filter_delay_line_delay_chain_4_n83,
         my_filter_delay_line_delay_chain_4_n82,
         my_filter_delay_line_delay_chain_4_n81,
         my_filter_delay_line_delay_chain_4_n80,
         my_filter_delay_line_delay_chain_4_n79,
         my_filter_delay_line_delay_chain_4_n78,
         my_filter_delay_line_delay_chain_4_n77,
         my_filter_delay_line_delay_chain_4_n76,
         my_filter_delay_line_delay_chain_4_n75,
         my_filter_delay_line_delay_chain_4_n74,
         my_filter_delay_line_delay_chain_4_n73,
         my_filter_delay_line_delay_chain_4_n72,
         my_filter_delay_line_delay_chain_4_n71,
         my_filter_delay_line_delay_chain_4_n70,
         my_filter_delay_line_delay_chain_4_n69,
         my_filter_delay_line_delay_chain_4_n68,
         my_filter_delay_line_delay_chain_4_n67,
         my_filter_delay_line_delay_chain_4_n66,
         my_filter_delay_line_delay_chain_4_n65,
         my_filter_delay_line_delay_chain_4_n64,
         my_filter_delay_line_delay_chain_4_n63,
         my_filter_delay_line_delay_chain_4_n62,
         my_filter_delay_line_delay_chain_4_n61,
         my_filter_delay_line_delay_chain_4_n60,
         my_filter_delay_line_delay_chain_4_n59,
         my_filter_delay_line_delay_chain_4_n58,
         my_filter_delay_line_delay_chain_4_n57,
         my_filter_delay_line_delay_chain_4_n56,
         my_filter_delay_line_delay_chain_4_n55,
         my_filter_delay_line_delay_chain_4_n54,
         my_filter_delay_line_delay_chain_4_n53,
         my_filter_delay_line_delay_chain_4_n52,
         my_filter_delay_line_delay_chain_4_n51,
         my_filter_delay_line_delay_chain_4_n50,
         my_filter_delay_line_delay_chain_4_n49,
         my_filter_delay_line_delay_chain_4_n48,
         my_filter_delay_line_delay_chain_5_n94,
         my_filter_delay_line_delay_chain_5_n93,
         my_filter_delay_line_delay_chain_5_n92,
         my_filter_delay_line_delay_chain_5_n91,
         my_filter_delay_line_delay_chain_5_n90,
         my_filter_delay_line_delay_chain_5_n89,
         my_filter_delay_line_delay_chain_5_n88,
         my_filter_delay_line_delay_chain_5_n87,
         my_filter_delay_line_delay_chain_5_n86,
         my_filter_delay_line_delay_chain_5_n85,
         my_filter_delay_line_delay_chain_5_n84,
         my_filter_delay_line_delay_chain_5_n83,
         my_filter_delay_line_delay_chain_5_n82,
         my_filter_delay_line_delay_chain_5_n81,
         my_filter_delay_line_delay_chain_5_n80,
         my_filter_delay_line_delay_chain_5_n79,
         my_filter_delay_line_delay_chain_5_n78,
         my_filter_delay_line_delay_chain_5_n77,
         my_filter_delay_line_delay_chain_5_n76,
         my_filter_delay_line_delay_chain_5_n75,
         my_filter_delay_line_delay_chain_5_n74,
         my_filter_delay_line_delay_chain_5_n73,
         my_filter_delay_line_delay_chain_5_n72,
         my_filter_delay_line_delay_chain_5_n71,
         my_filter_delay_line_delay_chain_5_n70,
         my_filter_delay_line_delay_chain_5_n69,
         my_filter_delay_line_delay_chain_5_n68,
         my_filter_delay_line_delay_chain_5_n67,
         my_filter_delay_line_delay_chain_5_n66,
         my_filter_delay_line_delay_chain_5_n65,
         my_filter_delay_line_delay_chain_5_n64,
         my_filter_delay_line_delay_chain_5_n63,
         my_filter_delay_line_delay_chain_5_n62,
         my_filter_delay_line_delay_chain_5_n61,
         my_filter_delay_line_delay_chain_5_n60,
         my_filter_delay_line_delay_chain_5_n59,
         my_filter_delay_line_delay_chain_5_n58,
         my_filter_delay_line_delay_chain_5_n57,
         my_filter_delay_line_delay_chain_5_n56,
         my_filter_delay_line_delay_chain_5_n55,
         my_filter_delay_line_delay_chain_5_n54,
         my_filter_delay_line_delay_chain_5_n53,
         my_filter_delay_line_delay_chain_5_n52,
         my_filter_delay_line_delay_chain_5_n51,
         my_filter_delay_line_delay_chain_5_n50,
         my_filter_delay_line_delay_chain_5_n49,
         my_filter_delay_line_delay_chain_5_n48,
         my_filter_delay_line_delay_chain_6_n93,
         my_filter_delay_line_delay_chain_6_n92,
         my_filter_delay_line_delay_chain_6_n91,
         my_filter_delay_line_delay_chain_6_n90,
         my_filter_delay_line_delay_chain_6_n89,
         my_filter_delay_line_delay_chain_6_n88,
         my_filter_delay_line_delay_chain_6_n87,
         my_filter_delay_line_delay_chain_6_n86,
         my_filter_delay_line_delay_chain_6_n85,
         my_filter_delay_line_delay_chain_6_n84,
         my_filter_delay_line_delay_chain_6_n83,
         my_filter_delay_line_delay_chain_6_n82,
         my_filter_delay_line_delay_chain_6_n81,
         my_filter_delay_line_delay_chain_6_n80,
         my_filter_delay_line_delay_chain_6_n79,
         my_filter_delay_line_delay_chain_6_n78,
         my_filter_delay_line_delay_chain_6_n77,
         my_filter_delay_line_delay_chain_6_n76,
         my_filter_delay_line_delay_chain_6_n75,
         my_filter_delay_line_delay_chain_6_n74,
         my_filter_delay_line_delay_chain_6_n73,
         my_filter_delay_line_delay_chain_6_n72,
         my_filter_delay_line_delay_chain_6_n71,
         my_filter_delay_line_delay_chain_6_n70,
         my_filter_delay_line_delay_chain_6_n69,
         my_filter_delay_line_delay_chain_6_n68,
         my_filter_delay_line_delay_chain_6_n67,
         my_filter_delay_line_delay_chain_6_n66,
         my_filter_delay_line_delay_chain_6_n65,
         my_filter_delay_line_delay_chain_6_n64,
         my_filter_delay_line_delay_chain_6_n63,
         my_filter_delay_line_delay_chain_6_n62,
         my_filter_delay_line_delay_chain_6_n61,
         my_filter_delay_line_delay_chain_6_n60,
         my_filter_delay_line_delay_chain_6_n59,
         my_filter_delay_line_delay_chain_6_n58,
         my_filter_delay_line_delay_chain_6_n57,
         my_filter_delay_line_delay_chain_6_n56,
         my_filter_delay_line_delay_chain_6_n55,
         my_filter_delay_line_delay_chain_6_n54,
         my_filter_delay_line_delay_chain_6_n53,
         my_filter_delay_line_delay_chain_6_n52,
         my_filter_delay_line_delay_chain_6_n51,
         my_filter_delay_line_delay_chain_6_n50,
         my_filter_delay_line_delay_chain_6_n49,
         my_filter_delay_line_delay_chain_6_n48,
         my_filter_delay_line_delay_chain_7_n93,
         my_filter_delay_line_delay_chain_7_n92,
         my_filter_delay_line_delay_chain_7_n91,
         my_filter_delay_line_delay_chain_7_n90,
         my_filter_delay_line_delay_chain_7_n89,
         my_filter_delay_line_delay_chain_7_n88,
         my_filter_delay_line_delay_chain_7_n87,
         my_filter_delay_line_delay_chain_7_n86,
         my_filter_delay_line_delay_chain_7_n85,
         my_filter_delay_line_delay_chain_7_n84,
         my_filter_delay_line_delay_chain_7_n83,
         my_filter_delay_line_delay_chain_7_n82,
         my_filter_delay_line_delay_chain_7_n81,
         my_filter_delay_line_delay_chain_7_n80,
         my_filter_delay_line_delay_chain_7_n79,
         my_filter_delay_line_delay_chain_7_n78,
         my_filter_delay_line_delay_chain_7_n77,
         my_filter_delay_line_delay_chain_7_n76,
         my_filter_delay_line_delay_chain_7_n75,
         my_filter_delay_line_delay_chain_7_n74,
         my_filter_delay_line_delay_chain_7_n73,
         my_filter_delay_line_delay_chain_7_n72,
         my_filter_delay_line_delay_chain_7_n71,
         my_filter_delay_line_delay_chain_7_n70,
         my_filter_delay_line_delay_chain_7_n69,
         my_filter_delay_line_delay_chain_7_n68,
         my_filter_delay_line_delay_chain_7_n67,
         my_filter_delay_line_delay_chain_7_n66,
         my_filter_delay_line_delay_chain_7_n65,
         my_filter_delay_line_delay_chain_7_n64,
         my_filter_delay_line_delay_chain_7_n63,
         my_filter_delay_line_delay_chain_7_n62,
         my_filter_delay_line_delay_chain_7_n61,
         my_filter_delay_line_delay_chain_7_n60,
         my_filter_delay_line_delay_chain_7_n59,
         my_filter_delay_line_delay_chain_7_n58,
         my_filter_delay_line_delay_chain_7_n57,
         my_filter_delay_line_delay_chain_7_n56,
         my_filter_delay_line_delay_chain_7_n55,
         my_filter_delay_line_delay_chain_7_n54,
         my_filter_delay_line_delay_chain_7_n53,
         my_filter_delay_line_delay_chain_7_n52,
         my_filter_delay_line_delay_chain_7_n51,
         my_filter_delay_line_delay_chain_7_n50,
         my_filter_delay_line_delay_chain_7_n49,
         my_filter_delay_line_delay_chain_7_n48,
         my_filter_delay_line_delay_chain_8_n93,
         my_filter_delay_line_delay_chain_8_n92,
         my_filter_delay_line_delay_chain_8_n91,
         my_filter_delay_line_delay_chain_8_n90,
         my_filter_delay_line_delay_chain_8_n89,
         my_filter_delay_line_delay_chain_8_n88,
         my_filter_delay_line_delay_chain_8_n87,
         my_filter_delay_line_delay_chain_8_n86,
         my_filter_delay_line_delay_chain_8_n85,
         my_filter_delay_line_delay_chain_8_n84,
         my_filter_delay_line_delay_chain_8_n83,
         my_filter_delay_line_delay_chain_8_n82,
         my_filter_delay_line_delay_chain_8_n81,
         my_filter_delay_line_delay_chain_8_n80,
         my_filter_delay_line_delay_chain_8_n79,
         my_filter_delay_line_delay_chain_8_n78,
         my_filter_delay_line_delay_chain_8_n77,
         my_filter_delay_line_delay_chain_8_n76,
         my_filter_delay_line_delay_chain_8_n75,
         my_filter_delay_line_delay_chain_8_n74,
         my_filter_delay_line_delay_chain_8_n73,
         my_filter_delay_line_delay_chain_8_n72,
         my_filter_delay_line_delay_chain_8_n71,
         my_filter_delay_line_delay_chain_8_n70,
         my_filter_delay_line_delay_chain_8_n69,
         my_filter_delay_line_delay_chain_8_n68,
         my_filter_delay_line_delay_chain_8_n67,
         my_filter_delay_line_delay_chain_8_n66,
         my_filter_delay_line_delay_chain_8_n65,
         my_filter_delay_line_delay_chain_8_n64,
         my_filter_delay_line_delay_chain_8_n63,
         my_filter_delay_line_delay_chain_8_n62,
         my_filter_delay_line_delay_chain_8_n61,
         my_filter_delay_line_delay_chain_8_n60,
         my_filter_delay_line_delay_chain_8_n59,
         my_filter_delay_line_delay_chain_8_n58,
         my_filter_delay_line_delay_chain_8_n57,
         my_filter_delay_line_delay_chain_8_n56,
         my_filter_delay_line_delay_chain_8_n55,
         my_filter_delay_line_delay_chain_8_n54,
         my_filter_delay_line_delay_chain_8_n53,
         my_filter_delay_line_delay_chain_8_n52,
         my_filter_delay_line_delay_chain_8_n51,
         my_filter_delay_line_delay_chain_8_n50,
         my_filter_delay_line_delay_chain_8_n49,
         my_filter_delay_line_delay_chain_8_n48,
         my_filter_delay_line_delay_chain_9_n93,
         my_filter_delay_line_delay_chain_9_n92,
         my_filter_delay_line_delay_chain_9_n91,
         my_filter_delay_line_delay_chain_9_n90,
         my_filter_delay_line_delay_chain_9_n89,
         my_filter_delay_line_delay_chain_9_n88,
         my_filter_delay_line_delay_chain_9_n87,
         my_filter_delay_line_delay_chain_9_n86,
         my_filter_delay_line_delay_chain_9_n85,
         my_filter_delay_line_delay_chain_9_n84,
         my_filter_delay_line_delay_chain_9_n83,
         my_filter_delay_line_delay_chain_9_n82,
         my_filter_delay_line_delay_chain_9_n81,
         my_filter_delay_line_delay_chain_9_n80,
         my_filter_delay_line_delay_chain_9_n79,
         my_filter_delay_line_delay_chain_9_n78,
         my_filter_delay_line_delay_chain_9_n77,
         my_filter_delay_line_delay_chain_9_n76,
         my_filter_delay_line_delay_chain_9_n75,
         my_filter_delay_line_delay_chain_9_n74,
         my_filter_delay_line_delay_chain_9_n73,
         my_filter_delay_line_delay_chain_9_n72,
         my_filter_delay_line_delay_chain_9_n71,
         my_filter_delay_line_delay_chain_9_n70,
         my_filter_delay_line_delay_chain_9_n69,
         my_filter_delay_line_delay_chain_9_n68,
         my_filter_delay_line_delay_chain_9_n67,
         my_filter_delay_line_delay_chain_9_n66,
         my_filter_delay_line_delay_chain_9_n65,
         my_filter_delay_line_delay_chain_9_n64,
         my_filter_delay_line_delay_chain_9_n63,
         my_filter_delay_line_delay_chain_9_n62,
         my_filter_delay_line_delay_chain_9_n61,
         my_filter_delay_line_delay_chain_9_n60,
         my_filter_delay_line_delay_chain_9_n59,
         my_filter_delay_line_delay_chain_9_n58,
         my_filter_delay_line_delay_chain_9_n57,
         my_filter_delay_line_delay_chain_9_n56,
         my_filter_delay_line_delay_chain_9_n55,
         my_filter_delay_line_delay_chain_9_n54,
         my_filter_delay_line_delay_chain_9_n53,
         my_filter_delay_line_delay_chain_9_n52,
         my_filter_delay_line_delay_chain_9_n51,
         my_filter_delay_line_delay_chain_9_n50,
         my_filter_delay_line_delay_chain_9_n49,
         my_filter_delay_line_delay_chain_9_n48,
         my_filter_first_coeff_mult_21_n113,
         my_filter_first_coeff_mult_21_n112,
         my_filter_first_coeff_mult_21_n111,
         my_filter_first_coeff_mult_21_n110,
         my_filter_first_coeff_mult_21_n109,
         my_filter_first_coeff_mult_21_n108,
         my_filter_first_coeff_mult_21_n107,
         my_filter_first_coeff_mult_21_n106,
         my_filter_first_coeff_mult_21_n105,
         my_filter_first_coeff_mult_21_n104,
         my_filter_first_coeff_mult_21_n103,
         my_filter_first_coeff_mult_21_n102,
         my_filter_first_coeff_mult_21_n101,
         my_filter_first_coeff_mult_21_n100, my_filter_first_coeff_mult_21_n99,
         my_filter_first_coeff_mult_21_n98, my_filter_first_coeff_mult_21_n97,
         my_filter_first_coeff_mult_21_n96, my_filter_first_coeff_mult_21_n95,
         my_filter_first_coeff_mult_21_n94, my_filter_first_coeff_mult_21_n93,
         my_filter_first_coeff_mult_21_n92, my_filter_first_coeff_mult_21_n91,
         my_filter_first_coeff_mult_21_n90, my_filter_first_coeff_mult_21_n89,
         my_filter_first_coeff_mult_21_n88, my_filter_first_coeff_mult_21_n87,
         my_filter_first_coeff_mult_21_n86, my_filter_first_coeff_mult_21_n85,
         my_filter_first_coeff_mult_21_n52, my_filter_first_coeff_mult_21_n51,
         my_filter_first_coeff_mult_21_n50, my_filter_first_coeff_mult_21_n49,
         my_filter_first_coeff_mult_21_n48, my_filter_first_coeff_mult_21_n47,
         my_filter_first_coeff_mult_21_n46, my_filter_first_coeff_mult_21_n45,
         my_filter_first_coeff_mult_21_n44, my_filter_first_coeff_mult_21_n43,
         my_filter_first_coeff_mult_21_n42, my_filter_first_coeff_mult_21_n41,
         my_filter_first_coeff_mult_21_n40, my_filter_first_coeff_mult_21_n39,
         my_filter_first_coeff_mult_21_n38, my_filter_first_coeff_mult_21_n37,
         my_filter_first_coeff_mult_21_n36, my_filter_first_coeff_mult_21_n35,
         my_filter_first_coeff_mult_21_n34, my_filter_first_coeff_mult_21_n33,
         my_filter_first_coeff_mult_21_n32, my_filter_first_coeff_mult_21_n31,
         my_filter_first_coeff_mult_21_n30, my_filter_first_coeff_mult_21_n29,
         my_filter_first_coeff_mult_21_n28, my_filter_first_coeff_mult_21_n27,
         my_filter_first_coeff_mult_21_n26, my_filter_first_coeff_mult_21_n25,
         my_filter_first_coeff_mult_21_n24, my_filter_first_coeff_mult_21_n23,
         my_filter_first_coeff_mult_21_n22, my_filter_first_coeff_mult_21_n21,
         my_filter_first_coeff_mult_21_n20, my_filter_first_coeff_mult_21_n19,
         my_filter_first_coeff_mult_21_n18, my_filter_first_coeff_mult_21_n17,
         my_filter_first_coeff_mult_21_n16, my_filter_first_coeff_mult_21_n15,
         my_filter_first_coeff_mult_21_n14, my_filter_first_coeff_mult_21_n13,
         my_filter_first_coeff_mult_21_n12, my_filter_first_coeff_mult_21_n11,
         my_filter_first_coeff_mult_21_n10, my_filter_first_coeff_mult_21_n9,
         my_filter_first_coeff_mult_21_n8, my_filter_first_coeff_mult_21_n7,
         my_filter_first_coeff_mult_21_n6, my_filter_first_coeff_mult_21_n5,
         my_filter_first_coeff_mult_21_n4, my_filter_first_coeff_mult_21_n3,
         my_filter_first_coeff_mult_21_A2_12_,
         my_filter_first_coeff_mult_21_A1_0_,
         my_filter_first_coeff_mult_21_A1_1_,
         my_filter_first_coeff_mult_21_A1_2_,
         my_filter_first_coeff_mult_21_A1_3_,
         my_filter_first_coeff_mult_21_A1_4_,
         my_filter_first_coeff_mult_21_A1_5_,
         my_filter_first_coeff_mult_21_A1_6_,
         my_filter_first_coeff_mult_21_A1_7_,
         my_filter_first_coeff_mult_21_A1_8_,
         my_filter_first_coeff_mult_21_A1_9_,
         my_filter_first_coeff_mult_21_A1_10_,
         my_filter_first_coeff_mult_21_SUMB_2__1_,
         my_filter_first_coeff_mult_21_SUMB_2__2_,
         my_filter_first_coeff_mult_21_SUMB_2__3_,
         my_filter_first_coeff_mult_21_SUMB_2__4_,
         my_filter_first_coeff_mult_21_SUMB_2__5_,
         my_filter_first_coeff_mult_21_SUMB_2__6_,
         my_filter_first_coeff_mult_21_SUMB_2__7_,
         my_filter_first_coeff_mult_21_SUMB_2__8_,
         my_filter_first_coeff_mult_21_SUMB_2__9_,
         my_filter_first_coeff_mult_21_SUMB_2__10_,
         my_filter_first_coeff_mult_21_SUMB_2__11_,
         my_filter_first_coeff_mult_21_SUMB_2__12_,
         my_filter_first_coeff_mult_21_SUMB_3__1_,
         my_filter_first_coeff_mult_21_SUMB_3__2_,
         my_filter_first_coeff_mult_21_SUMB_3__3_,
         my_filter_first_coeff_mult_21_SUMB_3__4_,
         my_filter_first_coeff_mult_21_SUMB_3__5_,
         my_filter_first_coeff_mult_21_SUMB_3__6_,
         my_filter_first_coeff_mult_21_SUMB_3__7_,
         my_filter_first_coeff_mult_21_SUMB_3__8_,
         my_filter_first_coeff_mult_21_SUMB_3__9_,
         my_filter_first_coeff_mult_21_SUMB_3__10_,
         my_filter_first_coeff_mult_21_SUMB_3__11_,
         my_filter_first_coeff_mult_21_SUMB_3__12_,
         my_filter_first_coeff_mult_21_SUMB_4__1_,
         my_filter_first_coeff_mult_21_SUMB_4__2_,
         my_filter_first_coeff_mult_21_SUMB_4__3_,
         my_filter_first_coeff_mult_21_SUMB_4__4_,
         my_filter_first_coeff_mult_21_SUMB_4__5_,
         my_filter_first_coeff_mult_21_SUMB_4__6_,
         my_filter_first_coeff_mult_21_SUMB_4__7_,
         my_filter_first_coeff_mult_21_SUMB_4__8_,
         my_filter_first_coeff_mult_21_SUMB_4__9_,
         my_filter_first_coeff_mult_21_SUMB_4__10_,
         my_filter_first_coeff_mult_21_SUMB_4__11_,
         my_filter_first_coeff_mult_21_SUMB_4__12_,
         my_filter_first_coeff_mult_21_SUMB_5__1_,
         my_filter_first_coeff_mult_21_SUMB_5__2_,
         my_filter_first_coeff_mult_21_SUMB_5__3_,
         my_filter_first_coeff_mult_21_SUMB_5__4_,
         my_filter_first_coeff_mult_21_SUMB_5__5_,
         my_filter_first_coeff_mult_21_SUMB_5__6_,
         my_filter_first_coeff_mult_21_SUMB_5__7_,
         my_filter_first_coeff_mult_21_SUMB_5__8_,
         my_filter_first_coeff_mult_21_SUMB_5__9_,
         my_filter_first_coeff_mult_21_SUMB_5__10_,
         my_filter_first_coeff_mult_21_SUMB_5__11_,
         my_filter_first_coeff_mult_21_SUMB_5__12_,
         my_filter_first_coeff_mult_21_SUMB_6__1_,
         my_filter_first_coeff_mult_21_SUMB_6__2_,
         my_filter_first_coeff_mult_21_SUMB_6__3_,
         my_filter_first_coeff_mult_21_SUMB_6__4_,
         my_filter_first_coeff_mult_21_SUMB_6__5_,
         my_filter_first_coeff_mult_21_SUMB_6__6_,
         my_filter_first_coeff_mult_21_SUMB_6__7_,
         my_filter_first_coeff_mult_21_SUMB_6__8_,
         my_filter_first_coeff_mult_21_SUMB_6__9_,
         my_filter_first_coeff_mult_21_SUMB_6__10_,
         my_filter_first_coeff_mult_21_SUMB_6__11_,
         my_filter_first_coeff_mult_21_SUMB_6__12_,
         my_filter_first_coeff_mult_21_SUMB_7__1_,
         my_filter_first_coeff_mult_21_SUMB_7__2_,
         my_filter_first_coeff_mult_21_SUMB_7__3_,
         my_filter_first_coeff_mult_21_SUMB_7__4_,
         my_filter_first_coeff_mult_21_SUMB_7__5_,
         my_filter_first_coeff_mult_21_SUMB_7__6_,
         my_filter_first_coeff_mult_21_SUMB_7__7_,
         my_filter_first_coeff_mult_21_SUMB_7__8_,
         my_filter_first_coeff_mult_21_SUMB_7__9_,
         my_filter_first_coeff_mult_21_SUMB_7__10_,
         my_filter_first_coeff_mult_21_SUMB_7__11_,
         my_filter_first_coeff_mult_21_SUMB_7__12_,
         my_filter_first_coeff_mult_21_SUMB_8__1_,
         my_filter_first_coeff_mult_21_SUMB_8__2_,
         my_filter_first_coeff_mult_21_SUMB_8__3_,
         my_filter_first_coeff_mult_21_SUMB_8__4_,
         my_filter_first_coeff_mult_21_SUMB_8__5_,
         my_filter_first_coeff_mult_21_SUMB_8__6_,
         my_filter_first_coeff_mult_21_SUMB_8__7_,
         my_filter_first_coeff_mult_21_SUMB_8__8_,
         my_filter_first_coeff_mult_21_SUMB_8__9_,
         my_filter_first_coeff_mult_21_SUMB_8__10_,
         my_filter_first_coeff_mult_21_SUMB_8__11_,
         my_filter_first_coeff_mult_21_SUMB_8__12_,
         my_filter_first_coeff_mult_21_SUMB_9__1_,
         my_filter_first_coeff_mult_21_SUMB_9__2_,
         my_filter_first_coeff_mult_21_SUMB_9__3_,
         my_filter_first_coeff_mult_21_SUMB_9__4_,
         my_filter_first_coeff_mult_21_SUMB_9__5_,
         my_filter_first_coeff_mult_21_SUMB_9__6_,
         my_filter_first_coeff_mult_21_SUMB_9__7_,
         my_filter_first_coeff_mult_21_SUMB_9__8_,
         my_filter_first_coeff_mult_21_SUMB_9__9_,
         my_filter_first_coeff_mult_21_SUMB_9__10_,
         my_filter_first_coeff_mult_21_SUMB_9__11_,
         my_filter_first_coeff_mult_21_SUMB_9__12_,
         my_filter_first_coeff_mult_21_SUMB_10__1_,
         my_filter_first_coeff_mult_21_SUMB_10__2_,
         my_filter_first_coeff_mult_21_SUMB_10__3_,
         my_filter_first_coeff_mult_21_SUMB_10__4_,
         my_filter_first_coeff_mult_21_SUMB_10__5_,
         my_filter_first_coeff_mult_21_SUMB_10__6_,
         my_filter_first_coeff_mult_21_SUMB_10__7_,
         my_filter_first_coeff_mult_21_SUMB_10__8_,
         my_filter_first_coeff_mult_21_SUMB_10__9_,
         my_filter_first_coeff_mult_21_SUMB_10__10_,
         my_filter_first_coeff_mult_21_SUMB_10__11_,
         my_filter_first_coeff_mult_21_SUMB_10__12_,
         my_filter_first_coeff_mult_21_SUMB_11__1_,
         my_filter_first_coeff_mult_21_SUMB_11__2_,
         my_filter_first_coeff_mult_21_SUMB_11__3_,
         my_filter_first_coeff_mult_21_SUMB_11__4_,
         my_filter_first_coeff_mult_21_SUMB_11__5_,
         my_filter_first_coeff_mult_21_SUMB_11__6_,
         my_filter_first_coeff_mult_21_SUMB_11__7_,
         my_filter_first_coeff_mult_21_SUMB_11__8_,
         my_filter_first_coeff_mult_21_SUMB_11__9_,
         my_filter_first_coeff_mult_21_SUMB_11__10_,
         my_filter_first_coeff_mult_21_SUMB_11__11_,
         my_filter_first_coeff_mult_21_SUMB_11__12_,
         my_filter_first_coeff_mult_21_SUMB_12__1_,
         my_filter_first_coeff_mult_21_SUMB_12__2_,
         my_filter_first_coeff_mult_21_SUMB_12__3_,
         my_filter_first_coeff_mult_21_SUMB_12__4_,
         my_filter_first_coeff_mult_21_SUMB_12__5_,
         my_filter_first_coeff_mult_21_SUMB_12__6_,
         my_filter_first_coeff_mult_21_SUMB_12__7_,
         my_filter_first_coeff_mult_21_SUMB_12__8_,
         my_filter_first_coeff_mult_21_SUMB_12__9_,
         my_filter_first_coeff_mult_21_SUMB_12__10_,
         my_filter_first_coeff_mult_21_SUMB_12__11_,
         my_filter_first_coeff_mult_21_SUMB_12__12_,
         my_filter_first_coeff_mult_21_SUMB_13__0_,
         my_filter_first_coeff_mult_21_SUMB_13__1_,
         my_filter_first_coeff_mult_21_SUMB_13__2_,
         my_filter_first_coeff_mult_21_SUMB_13__3_,
         my_filter_first_coeff_mult_21_SUMB_13__4_,
         my_filter_first_coeff_mult_21_SUMB_13__5_,
         my_filter_first_coeff_mult_21_SUMB_13__6_,
         my_filter_first_coeff_mult_21_SUMB_13__7_,
         my_filter_first_coeff_mult_21_SUMB_13__8_,
         my_filter_first_coeff_mult_21_SUMB_13__9_,
         my_filter_first_coeff_mult_21_SUMB_13__10_,
         my_filter_first_coeff_mult_21_SUMB_13__11_,
         my_filter_first_coeff_mult_21_SUMB_13__12_,
         my_filter_first_coeff_mult_21_SUMB_13__13_,
         my_filter_first_coeff_mult_21_CARRYB_1__0_,
         my_filter_first_coeff_mult_21_CARRYB_2__0_,
         my_filter_first_coeff_mult_21_CARRYB_2__1_,
         my_filter_first_coeff_mult_21_CARRYB_2__2_,
         my_filter_first_coeff_mult_21_CARRYB_2__3_,
         my_filter_first_coeff_mult_21_CARRYB_2__4_,
         my_filter_first_coeff_mult_21_CARRYB_2__5_,
         my_filter_first_coeff_mult_21_CARRYB_2__6_,
         my_filter_first_coeff_mult_21_CARRYB_2__7_,
         my_filter_first_coeff_mult_21_CARRYB_2__8_,
         my_filter_first_coeff_mult_21_CARRYB_2__9_,
         my_filter_first_coeff_mult_21_CARRYB_2__10_,
         my_filter_first_coeff_mult_21_CARRYB_2__11_,
         my_filter_first_coeff_mult_21_CARRYB_2__12_,
         my_filter_first_coeff_mult_21_CARRYB_3__0_,
         my_filter_first_coeff_mult_21_CARRYB_3__1_,
         my_filter_first_coeff_mult_21_CARRYB_3__2_,
         my_filter_first_coeff_mult_21_CARRYB_3__3_,
         my_filter_first_coeff_mult_21_CARRYB_3__4_,
         my_filter_first_coeff_mult_21_CARRYB_3__5_,
         my_filter_first_coeff_mult_21_CARRYB_3__6_,
         my_filter_first_coeff_mult_21_CARRYB_3__7_,
         my_filter_first_coeff_mult_21_CARRYB_3__8_,
         my_filter_first_coeff_mult_21_CARRYB_3__9_,
         my_filter_first_coeff_mult_21_CARRYB_3__10_,
         my_filter_first_coeff_mult_21_CARRYB_3__11_,
         my_filter_first_coeff_mult_21_CARRYB_3__12_,
         my_filter_first_coeff_mult_21_CARRYB_4__0_,
         my_filter_first_coeff_mult_21_CARRYB_4__1_,
         my_filter_first_coeff_mult_21_CARRYB_4__2_,
         my_filter_first_coeff_mult_21_CARRYB_4__3_,
         my_filter_first_coeff_mult_21_CARRYB_4__4_,
         my_filter_first_coeff_mult_21_CARRYB_4__5_,
         my_filter_first_coeff_mult_21_CARRYB_4__6_,
         my_filter_first_coeff_mult_21_CARRYB_4__7_,
         my_filter_first_coeff_mult_21_CARRYB_4__8_,
         my_filter_first_coeff_mult_21_CARRYB_4__9_,
         my_filter_first_coeff_mult_21_CARRYB_4__10_,
         my_filter_first_coeff_mult_21_CARRYB_4__11_,
         my_filter_first_coeff_mult_21_CARRYB_4__12_,
         my_filter_first_coeff_mult_21_CARRYB_5__0_,
         my_filter_first_coeff_mult_21_CARRYB_5__1_,
         my_filter_first_coeff_mult_21_CARRYB_5__2_,
         my_filter_first_coeff_mult_21_CARRYB_5__3_,
         my_filter_first_coeff_mult_21_CARRYB_5__4_,
         my_filter_first_coeff_mult_21_CARRYB_5__5_,
         my_filter_first_coeff_mult_21_CARRYB_5__6_,
         my_filter_first_coeff_mult_21_CARRYB_5__7_,
         my_filter_first_coeff_mult_21_CARRYB_5__8_,
         my_filter_first_coeff_mult_21_CARRYB_5__9_,
         my_filter_first_coeff_mult_21_CARRYB_5__10_,
         my_filter_first_coeff_mult_21_CARRYB_5__11_,
         my_filter_first_coeff_mult_21_CARRYB_5__12_,
         my_filter_first_coeff_mult_21_CARRYB_6__0_,
         my_filter_first_coeff_mult_21_CARRYB_6__1_,
         my_filter_first_coeff_mult_21_CARRYB_6__2_,
         my_filter_first_coeff_mult_21_CARRYB_6__3_,
         my_filter_first_coeff_mult_21_CARRYB_6__4_,
         my_filter_first_coeff_mult_21_CARRYB_6__5_,
         my_filter_first_coeff_mult_21_CARRYB_6__6_,
         my_filter_first_coeff_mult_21_CARRYB_6__7_,
         my_filter_first_coeff_mult_21_CARRYB_6__8_,
         my_filter_first_coeff_mult_21_CARRYB_6__9_,
         my_filter_first_coeff_mult_21_CARRYB_6__10_,
         my_filter_first_coeff_mult_21_CARRYB_6__11_,
         my_filter_first_coeff_mult_21_CARRYB_6__12_,
         my_filter_first_coeff_mult_21_CARRYB_7__0_,
         my_filter_first_coeff_mult_21_CARRYB_7__1_,
         my_filter_first_coeff_mult_21_CARRYB_7__2_,
         my_filter_first_coeff_mult_21_CARRYB_7__3_,
         my_filter_first_coeff_mult_21_CARRYB_7__4_,
         my_filter_first_coeff_mult_21_CARRYB_7__5_,
         my_filter_first_coeff_mult_21_CARRYB_7__6_,
         my_filter_first_coeff_mult_21_CARRYB_7__7_,
         my_filter_first_coeff_mult_21_CARRYB_7__8_,
         my_filter_first_coeff_mult_21_CARRYB_7__9_,
         my_filter_first_coeff_mult_21_CARRYB_7__10_,
         my_filter_first_coeff_mult_21_CARRYB_7__11_,
         my_filter_first_coeff_mult_21_CARRYB_7__12_,
         my_filter_first_coeff_mult_21_CARRYB_8__0_,
         my_filter_first_coeff_mult_21_CARRYB_8__1_,
         my_filter_first_coeff_mult_21_CARRYB_8__2_,
         my_filter_first_coeff_mult_21_CARRYB_8__3_,
         my_filter_first_coeff_mult_21_CARRYB_8__4_,
         my_filter_first_coeff_mult_21_CARRYB_8__5_,
         my_filter_first_coeff_mult_21_CARRYB_8__6_,
         my_filter_first_coeff_mult_21_CARRYB_8__7_,
         my_filter_first_coeff_mult_21_CARRYB_8__8_,
         my_filter_first_coeff_mult_21_CARRYB_8__9_,
         my_filter_first_coeff_mult_21_CARRYB_8__10_,
         my_filter_first_coeff_mult_21_CARRYB_8__11_,
         my_filter_first_coeff_mult_21_CARRYB_8__12_,
         my_filter_first_coeff_mult_21_CARRYB_9__0_,
         my_filter_first_coeff_mult_21_CARRYB_9__1_,
         my_filter_first_coeff_mult_21_CARRYB_9__2_,
         my_filter_first_coeff_mult_21_CARRYB_9__3_,
         my_filter_first_coeff_mult_21_CARRYB_9__4_,
         my_filter_first_coeff_mult_21_CARRYB_9__5_,
         my_filter_first_coeff_mult_21_CARRYB_9__6_,
         my_filter_first_coeff_mult_21_CARRYB_9__7_,
         my_filter_first_coeff_mult_21_CARRYB_9__8_,
         my_filter_first_coeff_mult_21_CARRYB_9__9_,
         my_filter_first_coeff_mult_21_CARRYB_9__10_,
         my_filter_first_coeff_mult_21_CARRYB_9__11_,
         my_filter_first_coeff_mult_21_CARRYB_9__12_,
         my_filter_first_coeff_mult_21_CARRYB_10__0_,
         my_filter_first_coeff_mult_21_CARRYB_10__1_,
         my_filter_first_coeff_mult_21_CARRYB_10__2_,
         my_filter_first_coeff_mult_21_CARRYB_10__3_,
         my_filter_first_coeff_mult_21_CARRYB_10__4_,
         my_filter_first_coeff_mult_21_CARRYB_10__5_,
         my_filter_first_coeff_mult_21_CARRYB_10__6_,
         my_filter_first_coeff_mult_21_CARRYB_10__7_,
         my_filter_first_coeff_mult_21_CARRYB_10__8_,
         my_filter_first_coeff_mult_21_CARRYB_10__9_,
         my_filter_first_coeff_mult_21_CARRYB_10__10_,
         my_filter_first_coeff_mult_21_CARRYB_10__11_,
         my_filter_first_coeff_mult_21_CARRYB_10__12_,
         my_filter_first_coeff_mult_21_CARRYB_11__0_,
         my_filter_first_coeff_mult_21_CARRYB_11__1_,
         my_filter_first_coeff_mult_21_CARRYB_11__2_,
         my_filter_first_coeff_mult_21_CARRYB_11__3_,
         my_filter_first_coeff_mult_21_CARRYB_11__4_,
         my_filter_first_coeff_mult_21_CARRYB_11__5_,
         my_filter_first_coeff_mult_21_CARRYB_11__6_,
         my_filter_first_coeff_mult_21_CARRYB_11__7_,
         my_filter_first_coeff_mult_21_CARRYB_11__8_,
         my_filter_first_coeff_mult_21_CARRYB_11__9_,
         my_filter_first_coeff_mult_21_CARRYB_11__10_,
         my_filter_first_coeff_mult_21_CARRYB_11__11_,
         my_filter_first_coeff_mult_21_CARRYB_11__12_,
         my_filter_first_coeff_mult_21_CARRYB_12__0_,
         my_filter_first_coeff_mult_21_CARRYB_12__1_,
         my_filter_first_coeff_mult_21_CARRYB_12__2_,
         my_filter_first_coeff_mult_21_CARRYB_12__3_,
         my_filter_first_coeff_mult_21_CARRYB_12__4_,
         my_filter_first_coeff_mult_21_CARRYB_12__5_,
         my_filter_first_coeff_mult_21_CARRYB_12__6_,
         my_filter_first_coeff_mult_21_CARRYB_12__7_,
         my_filter_first_coeff_mult_21_CARRYB_12__8_,
         my_filter_first_coeff_mult_21_CARRYB_12__9_,
         my_filter_first_coeff_mult_21_CARRYB_12__10_,
         my_filter_first_coeff_mult_21_CARRYB_12__11_,
         my_filter_first_coeff_mult_21_CARRYB_12__12_,
         my_filter_first_coeff_mult_21_CARRYB_13__0_,
         my_filter_first_coeff_mult_21_CARRYB_13__1_,
         my_filter_first_coeff_mult_21_CARRYB_13__2_,
         my_filter_first_coeff_mult_21_CARRYB_13__3_,
         my_filter_first_coeff_mult_21_CARRYB_13__4_,
         my_filter_first_coeff_mult_21_CARRYB_13__5_,
         my_filter_first_coeff_mult_21_CARRYB_13__6_,
         my_filter_first_coeff_mult_21_CARRYB_13__7_,
         my_filter_first_coeff_mult_21_CARRYB_13__8_,
         my_filter_first_coeff_mult_21_CARRYB_13__9_,
         my_filter_first_coeff_mult_21_CARRYB_13__10_,
         my_filter_first_coeff_mult_21_CARRYB_13__11_,
         my_filter_first_coeff_mult_21_CARRYB_13__12_,
         my_filter_first_coeff_mult_21_CARRYB_13__13_,
         my_filter_first_coeff_mult_21_ab_0__2_,
         my_filter_first_coeff_mult_21_ab_0__3_,
         my_filter_first_coeff_mult_21_ab_0__4_,
         my_filter_first_coeff_mult_21_ab_0__5_,
         my_filter_first_coeff_mult_21_ab_0__6_,
         my_filter_first_coeff_mult_21_ab_0__7_,
         my_filter_first_coeff_mult_21_ab_0__8_,
         my_filter_first_coeff_mult_21_ab_0__9_,
         my_filter_first_coeff_mult_21_ab_0__10_,
         my_filter_first_coeff_mult_21_ab_0__11_,
         my_filter_first_coeff_mult_21_ab_0__12_,
         my_filter_first_coeff_mult_21_ab_0__13_,
         my_filter_first_coeff_mult_21_ab_1__1_,
         my_filter_first_coeff_mult_21_ab_1__2_,
         my_filter_first_coeff_mult_21_ab_1__3_,
         my_filter_first_coeff_mult_21_ab_1__4_,
         my_filter_first_coeff_mult_21_ab_1__5_,
         my_filter_first_coeff_mult_21_ab_1__6_,
         my_filter_first_coeff_mult_21_ab_1__7_,
         my_filter_first_coeff_mult_21_ab_1__8_,
         my_filter_first_coeff_mult_21_ab_1__9_,
         my_filter_first_coeff_mult_21_ab_1__10_,
         my_filter_first_coeff_mult_21_ab_1__11_,
         my_filter_first_coeff_mult_21_ab_1__12_,
         my_filter_first_coeff_mult_21_ab_1__13_,
         my_filter_first_coeff_mult_21_ab_2__0_,
         my_filter_first_coeff_mult_21_ab_2__1_,
         my_filter_first_coeff_mult_21_ab_2__2_,
         my_filter_first_coeff_mult_21_ab_2__3_,
         my_filter_first_coeff_mult_21_ab_2__4_,
         my_filter_first_coeff_mult_21_ab_2__5_,
         my_filter_first_coeff_mult_21_ab_2__6_,
         my_filter_first_coeff_mult_21_ab_2__7_,
         my_filter_first_coeff_mult_21_ab_2__8_,
         my_filter_first_coeff_mult_21_ab_2__9_,
         my_filter_first_coeff_mult_21_ab_2__10_,
         my_filter_first_coeff_mult_21_ab_2__11_,
         my_filter_first_coeff_mult_21_ab_2__12_,
         my_filter_first_coeff_mult_21_ab_2__13_,
         my_filter_first_coeff_mult_21_ab_3__0_,
         my_filter_first_coeff_mult_21_ab_3__1_,
         my_filter_first_coeff_mult_21_ab_3__2_,
         my_filter_first_coeff_mult_21_ab_3__3_,
         my_filter_first_coeff_mult_21_ab_3__4_,
         my_filter_first_coeff_mult_21_ab_3__5_,
         my_filter_first_coeff_mult_21_ab_3__6_,
         my_filter_first_coeff_mult_21_ab_3__7_,
         my_filter_first_coeff_mult_21_ab_3__8_,
         my_filter_first_coeff_mult_21_ab_3__9_,
         my_filter_first_coeff_mult_21_ab_3__10_,
         my_filter_first_coeff_mult_21_ab_3__11_,
         my_filter_first_coeff_mult_21_ab_3__12_,
         my_filter_first_coeff_mult_21_ab_3__13_,
         my_filter_first_coeff_mult_21_ab_4__0_,
         my_filter_first_coeff_mult_21_ab_4__1_,
         my_filter_first_coeff_mult_21_ab_4__2_,
         my_filter_first_coeff_mult_21_ab_4__3_,
         my_filter_first_coeff_mult_21_ab_4__4_,
         my_filter_first_coeff_mult_21_ab_4__5_,
         my_filter_first_coeff_mult_21_ab_4__6_,
         my_filter_first_coeff_mult_21_ab_4__7_,
         my_filter_first_coeff_mult_21_ab_4__8_,
         my_filter_first_coeff_mult_21_ab_4__9_,
         my_filter_first_coeff_mult_21_ab_4__10_,
         my_filter_first_coeff_mult_21_ab_4__11_,
         my_filter_first_coeff_mult_21_ab_4__12_,
         my_filter_first_coeff_mult_21_ab_4__13_,
         my_filter_first_coeff_mult_21_ab_5__0_,
         my_filter_first_coeff_mult_21_ab_5__1_,
         my_filter_first_coeff_mult_21_ab_5__2_,
         my_filter_first_coeff_mult_21_ab_5__3_,
         my_filter_first_coeff_mult_21_ab_5__4_,
         my_filter_first_coeff_mult_21_ab_5__5_,
         my_filter_first_coeff_mult_21_ab_5__6_,
         my_filter_first_coeff_mult_21_ab_5__7_,
         my_filter_first_coeff_mult_21_ab_5__8_,
         my_filter_first_coeff_mult_21_ab_5__9_,
         my_filter_first_coeff_mult_21_ab_5__10_,
         my_filter_first_coeff_mult_21_ab_5__11_,
         my_filter_first_coeff_mult_21_ab_5__12_,
         my_filter_first_coeff_mult_21_ab_5__13_,
         my_filter_first_coeff_mult_21_ab_6__0_,
         my_filter_first_coeff_mult_21_ab_6__1_,
         my_filter_first_coeff_mult_21_ab_6__2_,
         my_filter_first_coeff_mult_21_ab_6__3_,
         my_filter_first_coeff_mult_21_ab_6__4_,
         my_filter_first_coeff_mult_21_ab_6__5_,
         my_filter_first_coeff_mult_21_ab_6__6_,
         my_filter_first_coeff_mult_21_ab_6__7_,
         my_filter_first_coeff_mult_21_ab_6__8_,
         my_filter_first_coeff_mult_21_ab_6__9_,
         my_filter_first_coeff_mult_21_ab_6__10_,
         my_filter_first_coeff_mult_21_ab_6__11_,
         my_filter_first_coeff_mult_21_ab_6__12_,
         my_filter_first_coeff_mult_21_ab_6__13_,
         my_filter_first_coeff_mult_21_ab_7__0_,
         my_filter_first_coeff_mult_21_ab_7__1_,
         my_filter_first_coeff_mult_21_ab_7__2_,
         my_filter_first_coeff_mult_21_ab_7__3_,
         my_filter_first_coeff_mult_21_ab_7__4_,
         my_filter_first_coeff_mult_21_ab_7__5_,
         my_filter_first_coeff_mult_21_ab_7__6_,
         my_filter_first_coeff_mult_21_ab_7__7_,
         my_filter_first_coeff_mult_21_ab_7__8_,
         my_filter_first_coeff_mult_21_ab_7__9_,
         my_filter_first_coeff_mult_21_ab_7__10_,
         my_filter_first_coeff_mult_21_ab_7__11_,
         my_filter_first_coeff_mult_21_ab_7__12_,
         my_filter_first_coeff_mult_21_ab_7__13_,
         my_filter_first_coeff_mult_21_ab_8__0_,
         my_filter_first_coeff_mult_21_ab_8__1_,
         my_filter_first_coeff_mult_21_ab_8__2_,
         my_filter_first_coeff_mult_21_ab_8__3_,
         my_filter_first_coeff_mult_21_ab_8__4_,
         my_filter_first_coeff_mult_21_ab_8__5_,
         my_filter_first_coeff_mult_21_ab_8__6_,
         my_filter_first_coeff_mult_21_ab_8__7_,
         my_filter_first_coeff_mult_21_ab_8__8_,
         my_filter_first_coeff_mult_21_ab_8__9_,
         my_filter_first_coeff_mult_21_ab_8__10_,
         my_filter_first_coeff_mult_21_ab_8__11_,
         my_filter_first_coeff_mult_21_ab_8__12_,
         my_filter_first_coeff_mult_21_ab_8__13_,
         my_filter_first_coeff_mult_21_ab_9__0_,
         my_filter_first_coeff_mult_21_ab_9__1_,
         my_filter_first_coeff_mult_21_ab_9__2_,
         my_filter_first_coeff_mult_21_ab_9__3_,
         my_filter_first_coeff_mult_21_ab_9__4_,
         my_filter_first_coeff_mult_21_ab_9__5_,
         my_filter_first_coeff_mult_21_ab_9__6_,
         my_filter_first_coeff_mult_21_ab_9__7_,
         my_filter_first_coeff_mult_21_ab_9__8_,
         my_filter_first_coeff_mult_21_ab_9__9_,
         my_filter_first_coeff_mult_21_ab_9__10_,
         my_filter_first_coeff_mult_21_ab_9__11_,
         my_filter_first_coeff_mult_21_ab_9__12_,
         my_filter_first_coeff_mult_21_ab_9__13_,
         my_filter_first_coeff_mult_21_ab_10__0_,
         my_filter_first_coeff_mult_21_ab_10__1_,
         my_filter_first_coeff_mult_21_ab_10__2_,
         my_filter_first_coeff_mult_21_ab_10__3_,
         my_filter_first_coeff_mult_21_ab_10__4_,
         my_filter_first_coeff_mult_21_ab_10__5_,
         my_filter_first_coeff_mult_21_ab_10__6_,
         my_filter_first_coeff_mult_21_ab_10__7_,
         my_filter_first_coeff_mult_21_ab_10__8_,
         my_filter_first_coeff_mult_21_ab_10__9_,
         my_filter_first_coeff_mult_21_ab_10__10_,
         my_filter_first_coeff_mult_21_ab_10__11_,
         my_filter_first_coeff_mult_21_ab_10__12_,
         my_filter_first_coeff_mult_21_ab_10__13_,
         my_filter_first_coeff_mult_21_ab_11__0_,
         my_filter_first_coeff_mult_21_ab_11__1_,
         my_filter_first_coeff_mult_21_ab_11__2_,
         my_filter_first_coeff_mult_21_ab_11__3_,
         my_filter_first_coeff_mult_21_ab_11__4_,
         my_filter_first_coeff_mult_21_ab_11__5_,
         my_filter_first_coeff_mult_21_ab_11__6_,
         my_filter_first_coeff_mult_21_ab_11__7_,
         my_filter_first_coeff_mult_21_ab_11__8_,
         my_filter_first_coeff_mult_21_ab_11__9_,
         my_filter_first_coeff_mult_21_ab_11__10_,
         my_filter_first_coeff_mult_21_ab_11__11_,
         my_filter_first_coeff_mult_21_ab_11__12_,
         my_filter_first_coeff_mult_21_ab_11__13_,
         my_filter_first_coeff_mult_21_ab_12__0_,
         my_filter_first_coeff_mult_21_ab_12__1_,
         my_filter_first_coeff_mult_21_ab_12__2_,
         my_filter_first_coeff_mult_21_ab_12__3_,
         my_filter_first_coeff_mult_21_ab_12__4_,
         my_filter_first_coeff_mult_21_ab_12__5_,
         my_filter_first_coeff_mult_21_ab_12__6_,
         my_filter_first_coeff_mult_21_ab_12__7_,
         my_filter_first_coeff_mult_21_ab_12__8_,
         my_filter_first_coeff_mult_21_ab_12__9_,
         my_filter_first_coeff_mult_21_ab_12__10_,
         my_filter_first_coeff_mult_21_ab_12__11_,
         my_filter_first_coeff_mult_21_ab_12__12_,
         my_filter_first_coeff_mult_21_ab_12__13_,
         my_filter_first_coeff_mult_21_ab_13__0_,
         my_filter_first_coeff_mult_21_ab_13__1_,
         my_filter_first_coeff_mult_21_ab_13__2_,
         my_filter_first_coeff_mult_21_ab_13__3_,
         my_filter_first_coeff_mult_21_ab_13__4_,
         my_filter_first_coeff_mult_21_ab_13__5_,
         my_filter_first_coeff_mult_21_ab_13__6_,
         my_filter_first_coeff_mult_21_ab_13__7_,
         my_filter_first_coeff_mult_21_ab_13__8_,
         my_filter_first_coeff_mult_21_ab_13__9_,
         my_filter_first_coeff_mult_21_ab_13__10_,
         my_filter_first_coeff_mult_21_ab_13__11_,
         my_filter_first_coeff_mult_21_ab_13__12_,
         my_filter_first_coeff_mult_21_ab_13__13_,
         my_filter_first_coeff_mult_21_FS_1_n70,
         my_filter_first_coeff_mult_21_FS_1_n69,
         my_filter_first_coeff_mult_21_FS_1_n68,
         my_filter_first_coeff_mult_21_FS_1_n67,
         my_filter_first_coeff_mult_21_FS_1_n66,
         my_filter_first_coeff_mult_21_FS_1_n65,
         my_filter_first_coeff_mult_21_FS_1_n64,
         my_filter_first_coeff_mult_21_FS_1_n63,
         my_filter_first_coeff_mult_21_FS_1_n62,
         my_filter_first_coeff_mult_21_FS_1_n61,
         my_filter_first_coeff_mult_21_FS_1_n60,
         my_filter_first_coeff_mult_21_FS_1_n59,
         my_filter_first_coeff_mult_21_FS_1_n58,
         my_filter_first_coeff_mult_21_FS_1_n57,
         my_filter_first_coeff_mult_21_FS_1_n56,
         my_filter_first_coeff_mult_21_FS_1_n55,
         my_filter_first_coeff_mult_21_FS_1_n54,
         my_filter_first_coeff_mult_21_FS_1_n53,
         my_filter_first_coeff_mult_21_FS_1_n52,
         my_filter_first_coeff_mult_21_FS_1_n51,
         my_filter_first_coeff_mult_21_FS_1_n50,
         my_filter_first_coeff_mult_21_FS_1_n49,
         my_filter_first_coeff_mult_21_FS_1_n48,
         my_filter_first_coeff_mult_21_FS_1_n47,
         my_filter_first_coeff_mult_21_FS_1_n46,
         my_filter_first_coeff_mult_21_FS_1_n45,
         my_filter_first_coeff_mult_21_FS_1_n44,
         my_filter_first_coeff_mult_21_FS_1_n43,
         my_filter_first_coeff_mult_21_FS_1_n42,
         my_filter_first_coeff_mult_21_FS_1_n41,
         my_filter_first_coeff_mult_21_FS_1_n40,
         my_filter_first_coeff_mult_21_FS_1_n39,
         my_filter_first_coeff_mult_21_FS_1_n38,
         my_filter_first_coeff_mult_21_FS_1_n37,
         my_filter_first_coeff_mult_21_FS_1_n36,
         my_filter_first_coeff_mult_21_FS_1_n35,
         my_filter_first_coeff_mult_21_FS_1_n34,
         my_filter_first_coeff_mult_21_FS_1_n33,
         my_filter_first_coeff_mult_21_FS_1_n32,
         my_filter_first_coeff_mult_21_FS_1_n31,
         my_filter_first_coeff_mult_21_FS_1_n30,
         my_filter_first_coeff_mult_21_FS_1_n29,
         my_filter_first_coeff_mult_21_FS_1_n28,
         my_filter_first_coeff_mult_21_FS_1_n27,
         my_filter_first_coeff_mult_21_FS_1_n26,
         my_filter_first_coeff_mult_21_FS_1_n25,
         my_filter_first_coeff_mult_21_FS_1_n24,
         my_filter_first_coeff_mult_21_FS_1_n23,
         my_filter_first_coeff_mult_21_FS_1_n22,
         my_filter_first_coeff_mult_21_FS_1_n21,
         my_filter_first_coeff_mult_21_FS_1_n20,
         my_filter_first_coeff_mult_21_FS_1_n19,
         my_filter_first_coeff_mult_21_FS_1_n18,
         my_filter_first_coeff_mult_21_FS_1_n17,
         my_filter_first_coeff_mult_21_FS_1_n16,
         my_filter_first_coeff_mult_21_FS_1_n15,
         my_filter_first_coeff_mult_21_FS_1_n14,
         my_filter_first_coeff_mult_21_FS_1_n13,
         my_filter_adder_mult_0_multiplication_mult_21_n113,
         my_filter_adder_mult_0_multiplication_mult_21_n112,
         my_filter_adder_mult_0_multiplication_mult_21_n111,
         my_filter_adder_mult_0_multiplication_mult_21_n110,
         my_filter_adder_mult_0_multiplication_mult_21_n109,
         my_filter_adder_mult_0_multiplication_mult_21_n108,
         my_filter_adder_mult_0_multiplication_mult_21_n107,
         my_filter_adder_mult_0_multiplication_mult_21_n106,
         my_filter_adder_mult_0_multiplication_mult_21_n105,
         my_filter_adder_mult_0_multiplication_mult_21_n104,
         my_filter_adder_mult_0_multiplication_mult_21_n103,
         my_filter_adder_mult_0_multiplication_mult_21_n102,
         my_filter_adder_mult_0_multiplication_mult_21_n101,
         my_filter_adder_mult_0_multiplication_mult_21_n100,
         my_filter_adder_mult_0_multiplication_mult_21_n99,
         my_filter_adder_mult_0_multiplication_mult_21_n98,
         my_filter_adder_mult_0_multiplication_mult_21_n97,
         my_filter_adder_mult_0_multiplication_mult_21_n96,
         my_filter_adder_mult_0_multiplication_mult_21_n95,
         my_filter_adder_mult_0_multiplication_mult_21_n94,
         my_filter_adder_mult_0_multiplication_mult_21_n93,
         my_filter_adder_mult_0_multiplication_mult_21_n92,
         my_filter_adder_mult_0_multiplication_mult_21_n91,
         my_filter_adder_mult_0_multiplication_mult_21_n90,
         my_filter_adder_mult_0_multiplication_mult_21_n89,
         my_filter_adder_mult_0_multiplication_mult_21_n88,
         my_filter_adder_mult_0_multiplication_mult_21_n87,
         my_filter_adder_mult_0_multiplication_mult_21_n86,
         my_filter_adder_mult_0_multiplication_mult_21_n85,
         my_filter_adder_mult_0_multiplication_mult_21_n52,
         my_filter_adder_mult_0_multiplication_mult_21_n51,
         my_filter_adder_mult_0_multiplication_mult_21_n50,
         my_filter_adder_mult_0_multiplication_mult_21_n49,
         my_filter_adder_mult_0_multiplication_mult_21_n48,
         my_filter_adder_mult_0_multiplication_mult_21_n47,
         my_filter_adder_mult_0_multiplication_mult_21_n46,
         my_filter_adder_mult_0_multiplication_mult_21_n45,
         my_filter_adder_mult_0_multiplication_mult_21_n44,
         my_filter_adder_mult_0_multiplication_mult_21_n43,
         my_filter_adder_mult_0_multiplication_mult_21_n42,
         my_filter_adder_mult_0_multiplication_mult_21_n41,
         my_filter_adder_mult_0_multiplication_mult_21_n40,
         my_filter_adder_mult_0_multiplication_mult_21_n39,
         my_filter_adder_mult_0_multiplication_mult_21_n38,
         my_filter_adder_mult_0_multiplication_mult_21_n37,
         my_filter_adder_mult_0_multiplication_mult_21_n36,
         my_filter_adder_mult_0_multiplication_mult_21_n35,
         my_filter_adder_mult_0_multiplication_mult_21_n34,
         my_filter_adder_mult_0_multiplication_mult_21_n33,
         my_filter_adder_mult_0_multiplication_mult_21_n32,
         my_filter_adder_mult_0_multiplication_mult_21_n31,
         my_filter_adder_mult_0_multiplication_mult_21_n30,
         my_filter_adder_mult_0_multiplication_mult_21_n29,
         my_filter_adder_mult_0_multiplication_mult_21_n28,
         my_filter_adder_mult_0_multiplication_mult_21_n27,
         my_filter_adder_mult_0_multiplication_mult_21_n26,
         my_filter_adder_mult_0_multiplication_mult_21_n25,
         my_filter_adder_mult_0_multiplication_mult_21_n24,
         my_filter_adder_mult_0_multiplication_mult_21_n23,
         my_filter_adder_mult_0_multiplication_mult_21_n22,
         my_filter_adder_mult_0_multiplication_mult_21_n21,
         my_filter_adder_mult_0_multiplication_mult_21_n20,
         my_filter_adder_mult_0_multiplication_mult_21_n19,
         my_filter_adder_mult_0_multiplication_mult_21_n18,
         my_filter_adder_mult_0_multiplication_mult_21_n17,
         my_filter_adder_mult_0_multiplication_mult_21_n16,
         my_filter_adder_mult_0_multiplication_mult_21_n15,
         my_filter_adder_mult_0_multiplication_mult_21_n14,
         my_filter_adder_mult_0_multiplication_mult_21_n13,
         my_filter_adder_mult_0_multiplication_mult_21_n12,
         my_filter_adder_mult_0_multiplication_mult_21_n11,
         my_filter_adder_mult_0_multiplication_mult_21_n10,
         my_filter_adder_mult_0_multiplication_mult_21_n9,
         my_filter_adder_mult_0_multiplication_mult_21_n8,
         my_filter_adder_mult_0_multiplication_mult_21_n7,
         my_filter_adder_mult_0_multiplication_mult_21_n6,
         my_filter_adder_mult_0_multiplication_mult_21_n5,
         my_filter_adder_mult_0_multiplication_mult_21_n4,
         my_filter_adder_mult_0_multiplication_mult_21_n3,
         my_filter_adder_mult_0_multiplication_mult_21_A2_12_,
         my_filter_adder_mult_0_multiplication_mult_21_A1_0_,
         my_filter_adder_mult_0_multiplication_mult_21_A1_1_,
         my_filter_adder_mult_0_multiplication_mult_21_A1_2_,
         my_filter_adder_mult_0_multiplication_mult_21_A1_3_,
         my_filter_adder_mult_0_multiplication_mult_21_A1_4_,
         my_filter_adder_mult_0_multiplication_mult_21_A1_5_,
         my_filter_adder_mult_0_multiplication_mult_21_A1_6_,
         my_filter_adder_mult_0_multiplication_mult_21_A1_7_,
         my_filter_adder_mult_0_multiplication_mult_21_A1_8_,
         my_filter_adder_mult_0_multiplication_mult_21_A1_9_,
         my_filter_adder_mult_0_multiplication_mult_21_A1_10_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_2__1_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_2__2_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_2__3_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_2__4_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_2__5_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_2__6_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_2__7_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_2__8_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_2__9_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_2__10_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_2__11_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_2__12_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_3__1_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_3__2_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_3__3_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_3__4_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_3__5_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_3__6_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_3__7_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_3__8_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_3__9_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_3__10_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_3__11_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_3__12_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_4__1_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_4__2_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_4__3_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_4__4_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_4__5_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_4__6_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_4__7_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_4__8_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_4__9_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_4__10_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_4__11_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_4__12_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_5__1_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_5__2_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_5__3_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_5__4_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_5__5_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_5__6_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_5__7_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_5__8_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_5__9_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_5__10_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_5__11_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_5__12_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_6__1_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_6__2_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_6__3_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_6__4_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_6__5_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_6__6_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_6__7_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_6__8_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_6__9_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_6__10_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_6__11_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_6__12_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_7__1_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_7__2_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_7__3_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_7__4_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_7__5_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_7__6_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_7__7_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_7__8_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_7__9_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_7__10_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_7__11_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_7__12_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_8__1_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_8__2_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_8__3_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_8__4_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_8__5_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_8__6_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_8__7_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_8__8_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_8__9_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_8__10_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_8__11_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_8__12_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_9__1_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_9__2_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_9__3_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_9__4_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_9__5_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_9__6_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_9__7_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_9__8_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_9__9_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_9__10_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_9__11_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_9__12_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_10__1_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_10__2_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_10__3_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_10__4_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_10__5_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_10__6_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_10__7_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_10__8_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_10__9_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_10__10_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_10__11_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_10__12_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_11__1_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_11__2_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_11__3_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_11__4_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_11__5_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_11__6_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_11__7_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_11__8_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_11__9_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_11__10_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_11__11_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_11__12_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_12__1_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_12__2_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_12__3_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_12__4_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_12__5_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_12__6_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_12__7_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_12__8_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_12__9_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_12__10_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_12__11_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_12__12_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_13__0_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_13__1_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_13__2_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_13__3_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_13__4_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_13__5_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_13__6_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_13__7_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_13__8_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_13__9_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_13__10_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_13__11_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_13__12_,
         my_filter_adder_mult_0_multiplication_mult_21_SUMB_13__13_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_1__0_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_2__0_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_2__1_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_2__2_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_2__3_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_2__4_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_2__5_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_2__6_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_2__7_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_2__8_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_2__9_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_2__10_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_2__11_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_2__12_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_3__0_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_3__1_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_3__2_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_3__3_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_3__4_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_3__5_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_3__6_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_3__7_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_3__8_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_3__9_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_3__10_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_3__11_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_3__12_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_4__0_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_4__1_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_4__2_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_4__3_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_4__4_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_4__5_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_4__6_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_4__7_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_4__8_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_4__9_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_4__10_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_4__11_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_4__12_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_5__0_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_5__1_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_5__2_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_5__3_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_5__4_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_5__5_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_5__6_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_5__7_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_5__8_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_5__9_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_5__10_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_5__11_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_5__12_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_6__0_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_6__1_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_6__2_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_6__3_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_6__4_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_6__5_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_6__6_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_6__7_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_6__8_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_6__9_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_6__10_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_6__11_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_6__12_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_7__0_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_7__1_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_7__2_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_7__3_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_7__4_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_7__5_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_7__6_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_7__7_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_7__8_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_7__9_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_7__10_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_7__11_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_7__12_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_8__0_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_8__1_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_8__2_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_8__3_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_8__4_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_8__5_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_8__6_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_8__7_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_8__8_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_8__9_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_8__10_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_8__11_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_8__12_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_9__0_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_9__1_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_9__2_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_9__3_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_9__4_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_9__5_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_9__6_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_9__7_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_9__8_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_9__9_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_9__10_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_9__11_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_9__12_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_10__0_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_10__1_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_10__2_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_10__3_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_10__4_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_10__5_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_10__6_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_10__7_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_10__8_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_10__9_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_10__10_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_10__11_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_10__12_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_11__0_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_11__1_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_11__2_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_11__3_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_11__4_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_11__5_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_11__6_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_11__7_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_11__8_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_11__9_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_11__10_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_11__11_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_11__12_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_12__0_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_12__1_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_12__2_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_12__3_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_12__4_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_12__5_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_12__6_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_12__7_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_12__8_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_12__9_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_12__10_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_12__11_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_12__12_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_13__0_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_13__1_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_13__2_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_13__3_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_13__4_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_13__5_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_13__6_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_13__7_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_13__8_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_13__9_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_13__10_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_13__11_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_13__12_,
         my_filter_adder_mult_0_multiplication_mult_21_CARRYB_13__13_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_0__2_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_0__3_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_0__4_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_0__5_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_0__6_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_0__7_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_0__8_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_0__9_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_0__10_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_0__11_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_0__12_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_0__13_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_1__1_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_1__2_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_1__3_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_1__4_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_1__5_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_1__6_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_1__7_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_1__8_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_1__9_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_1__10_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_1__11_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_1__12_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_1__13_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_2__0_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_2__1_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_2__2_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_2__3_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_2__4_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_2__5_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_2__6_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_2__7_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_2__8_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_2__9_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_2__10_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_2__11_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_2__12_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_2__13_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_3__0_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_3__1_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_3__2_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_3__3_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_3__4_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_3__5_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_3__6_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_3__7_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_3__8_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_3__9_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_3__10_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_3__11_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_3__12_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_3__13_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_4__0_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_4__1_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_4__2_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_4__3_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_4__4_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_4__5_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_4__6_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_4__7_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_4__8_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_4__9_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_4__10_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_4__11_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_4__12_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_4__13_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_5__0_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_5__1_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_5__2_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_5__3_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_5__4_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_5__5_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_5__6_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_5__7_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_5__8_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_5__9_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_5__10_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_5__11_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_5__12_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_5__13_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_6__0_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_6__1_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_6__2_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_6__3_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_6__4_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_6__5_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_6__6_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_6__7_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_6__8_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_6__9_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_6__10_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_6__11_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_6__12_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_6__13_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_7__0_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_7__1_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_7__2_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_7__3_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_7__4_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_7__5_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_7__6_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_7__7_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_7__8_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_7__9_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_7__10_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_7__11_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_7__12_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_7__13_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_8__0_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_8__1_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_8__2_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_8__3_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_8__4_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_8__5_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_8__6_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_8__7_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_8__8_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_8__9_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_8__10_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_8__11_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_8__12_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_8__13_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_9__0_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_9__1_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_9__2_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_9__3_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_9__4_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_9__5_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_9__6_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_9__7_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_9__8_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_9__9_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_9__10_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_9__11_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_9__12_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_9__13_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_10__0_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_10__1_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_10__2_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_10__3_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_10__4_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_10__5_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_10__6_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_10__7_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_10__8_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_10__9_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_10__10_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_10__11_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_10__12_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_10__13_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_11__0_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_11__1_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_11__2_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_11__3_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_11__4_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_11__5_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_11__6_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_11__7_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_11__8_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_11__9_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_11__10_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_11__11_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_11__12_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_11__13_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_12__0_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_12__1_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_12__2_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_12__3_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_12__4_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_12__5_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_12__6_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_12__7_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_12__8_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_12__9_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_12__10_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_12__11_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_12__12_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_12__13_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_13__0_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_13__1_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_13__2_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_13__3_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_13__4_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_13__5_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_13__6_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_13__7_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_13__8_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_13__9_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_13__10_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_13__11_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_13__12_,
         my_filter_adder_mult_0_multiplication_mult_21_ab_13__13_,
         my_filter_adder_mult_0_multiplication_mult_21_FS_1_n71,
         my_filter_adder_mult_0_multiplication_mult_21_FS_1_n70,
         my_filter_adder_mult_0_multiplication_mult_21_FS_1_n69,
         my_filter_adder_mult_0_multiplication_mult_21_FS_1_n68,
         my_filter_adder_mult_0_multiplication_mult_21_FS_1_n67,
         my_filter_adder_mult_0_multiplication_mult_21_FS_1_n66,
         my_filter_adder_mult_0_multiplication_mult_21_FS_1_n65,
         my_filter_adder_mult_0_multiplication_mult_21_FS_1_n64,
         my_filter_adder_mult_0_multiplication_mult_21_FS_1_n63,
         my_filter_adder_mult_0_multiplication_mult_21_FS_1_n62,
         my_filter_adder_mult_0_multiplication_mult_21_FS_1_n60,
         my_filter_adder_mult_0_multiplication_mult_21_FS_1_n59,
         my_filter_adder_mult_0_multiplication_mult_21_FS_1_n58,
         my_filter_adder_mult_0_multiplication_mult_21_FS_1_n57,
         my_filter_adder_mult_0_multiplication_mult_21_FS_1_n56,
         my_filter_adder_mult_0_multiplication_mult_21_FS_1_n55,
         my_filter_adder_mult_0_multiplication_mult_21_FS_1_n54,
         my_filter_adder_mult_0_multiplication_mult_21_FS_1_n53,
         my_filter_adder_mult_0_multiplication_mult_21_FS_1_n52,
         my_filter_adder_mult_0_multiplication_mult_21_FS_1_n51,
         my_filter_adder_mult_0_multiplication_mult_21_FS_1_n50,
         my_filter_adder_mult_0_multiplication_mult_21_FS_1_n49,
         my_filter_adder_mult_0_multiplication_mult_21_FS_1_n48,
         my_filter_adder_mult_0_multiplication_mult_21_FS_1_n47,
         my_filter_adder_mult_0_multiplication_mult_21_FS_1_n46,
         my_filter_adder_mult_0_multiplication_mult_21_FS_1_n45,
         my_filter_adder_mult_0_multiplication_mult_21_FS_1_n44,
         my_filter_adder_mult_0_multiplication_mult_21_FS_1_n43,
         my_filter_adder_mult_0_multiplication_mult_21_FS_1_n42,
         my_filter_adder_mult_0_multiplication_mult_21_FS_1_n41,
         my_filter_adder_mult_0_multiplication_mult_21_FS_1_n40,
         my_filter_adder_mult_0_multiplication_mult_21_FS_1_n39,
         my_filter_adder_mult_0_multiplication_mult_21_FS_1_n38,
         my_filter_adder_mult_0_multiplication_mult_21_FS_1_n37,
         my_filter_adder_mult_0_multiplication_mult_21_FS_1_n36,
         my_filter_adder_mult_0_multiplication_mult_21_FS_1_n35,
         my_filter_adder_mult_0_multiplication_mult_21_FS_1_n34,
         my_filter_adder_mult_0_multiplication_mult_21_FS_1_n33,
         my_filter_adder_mult_0_multiplication_mult_21_FS_1_n32,
         my_filter_adder_mult_0_multiplication_mult_21_FS_1_n31,
         my_filter_adder_mult_0_multiplication_mult_21_FS_1_n30,
         my_filter_adder_mult_0_multiplication_mult_21_FS_1_n29,
         my_filter_adder_mult_0_multiplication_mult_21_FS_1_n28,
         my_filter_adder_mult_0_multiplication_mult_21_FS_1_n27,
         my_filter_adder_mult_0_multiplication_mult_21_FS_1_n26,
         my_filter_adder_mult_0_multiplication_mult_21_FS_1_n25,
         my_filter_adder_mult_0_multiplication_mult_21_FS_1_n24,
         my_filter_adder_mult_0_multiplication_mult_21_FS_1_n23,
         my_filter_adder_mult_0_multiplication_mult_21_FS_1_n22,
         my_filter_adder_mult_0_multiplication_mult_21_FS_1_n21,
         my_filter_adder_mult_0_multiplication_mult_21_FS_1_n20,
         my_filter_adder_mult_0_multiplication_mult_21_FS_1_n19,
         my_filter_adder_mult_0_multiplication_mult_21_FS_1_n18,
         my_filter_adder_mult_0_multiplication_mult_21_FS_1_n17,
         my_filter_adder_mult_0_multiplication_mult_21_FS_1_n16,
         my_filter_adder_mult_0_multiplication_mult_21_FS_1_n15,
         my_filter_adder_mult_0_multiplication_mult_21_FS_1_n14,
         my_filter_adder_mult_0_multiplication_mult_21_FS_1_n13,
         my_filter_adder_mult_0_addition_add_19_n1,
         my_filter_adder_mult_1_multiplication_mult_21_n113,
         my_filter_adder_mult_1_multiplication_mult_21_n112,
         my_filter_adder_mult_1_multiplication_mult_21_n111,
         my_filter_adder_mult_1_multiplication_mult_21_n110,
         my_filter_adder_mult_1_multiplication_mult_21_n109,
         my_filter_adder_mult_1_multiplication_mult_21_n108,
         my_filter_adder_mult_1_multiplication_mult_21_n107,
         my_filter_adder_mult_1_multiplication_mult_21_n106,
         my_filter_adder_mult_1_multiplication_mult_21_n105,
         my_filter_adder_mult_1_multiplication_mult_21_n104,
         my_filter_adder_mult_1_multiplication_mult_21_n103,
         my_filter_adder_mult_1_multiplication_mult_21_n102,
         my_filter_adder_mult_1_multiplication_mult_21_n101,
         my_filter_adder_mult_1_multiplication_mult_21_n100,
         my_filter_adder_mult_1_multiplication_mult_21_n99,
         my_filter_adder_mult_1_multiplication_mult_21_n98,
         my_filter_adder_mult_1_multiplication_mult_21_n97,
         my_filter_adder_mult_1_multiplication_mult_21_n96,
         my_filter_adder_mult_1_multiplication_mult_21_n95,
         my_filter_adder_mult_1_multiplication_mult_21_n94,
         my_filter_adder_mult_1_multiplication_mult_21_n93,
         my_filter_adder_mult_1_multiplication_mult_21_n92,
         my_filter_adder_mult_1_multiplication_mult_21_n91,
         my_filter_adder_mult_1_multiplication_mult_21_n90,
         my_filter_adder_mult_1_multiplication_mult_21_n89,
         my_filter_adder_mult_1_multiplication_mult_21_n88,
         my_filter_adder_mult_1_multiplication_mult_21_n87,
         my_filter_adder_mult_1_multiplication_mult_21_n86,
         my_filter_adder_mult_1_multiplication_mult_21_n85,
         my_filter_adder_mult_1_multiplication_mult_21_n52,
         my_filter_adder_mult_1_multiplication_mult_21_n51,
         my_filter_adder_mult_1_multiplication_mult_21_n50,
         my_filter_adder_mult_1_multiplication_mult_21_n49,
         my_filter_adder_mult_1_multiplication_mult_21_n48,
         my_filter_adder_mult_1_multiplication_mult_21_n47,
         my_filter_adder_mult_1_multiplication_mult_21_n46,
         my_filter_adder_mult_1_multiplication_mult_21_n45,
         my_filter_adder_mult_1_multiplication_mult_21_n44,
         my_filter_adder_mult_1_multiplication_mult_21_n43,
         my_filter_adder_mult_1_multiplication_mult_21_n42,
         my_filter_adder_mult_1_multiplication_mult_21_n41,
         my_filter_adder_mult_1_multiplication_mult_21_n40,
         my_filter_adder_mult_1_multiplication_mult_21_n39,
         my_filter_adder_mult_1_multiplication_mult_21_n38,
         my_filter_adder_mult_1_multiplication_mult_21_n37,
         my_filter_adder_mult_1_multiplication_mult_21_n36,
         my_filter_adder_mult_1_multiplication_mult_21_n35,
         my_filter_adder_mult_1_multiplication_mult_21_n34,
         my_filter_adder_mult_1_multiplication_mult_21_n33,
         my_filter_adder_mult_1_multiplication_mult_21_n32,
         my_filter_adder_mult_1_multiplication_mult_21_n31,
         my_filter_adder_mult_1_multiplication_mult_21_n30,
         my_filter_adder_mult_1_multiplication_mult_21_n29,
         my_filter_adder_mult_1_multiplication_mult_21_n28,
         my_filter_adder_mult_1_multiplication_mult_21_n27,
         my_filter_adder_mult_1_multiplication_mult_21_n26,
         my_filter_adder_mult_1_multiplication_mult_21_n25,
         my_filter_adder_mult_1_multiplication_mult_21_n24,
         my_filter_adder_mult_1_multiplication_mult_21_n23,
         my_filter_adder_mult_1_multiplication_mult_21_n22,
         my_filter_adder_mult_1_multiplication_mult_21_n21,
         my_filter_adder_mult_1_multiplication_mult_21_n20,
         my_filter_adder_mult_1_multiplication_mult_21_n19,
         my_filter_adder_mult_1_multiplication_mult_21_n18,
         my_filter_adder_mult_1_multiplication_mult_21_n17,
         my_filter_adder_mult_1_multiplication_mult_21_n16,
         my_filter_adder_mult_1_multiplication_mult_21_n15,
         my_filter_adder_mult_1_multiplication_mult_21_n14,
         my_filter_adder_mult_1_multiplication_mult_21_n13,
         my_filter_adder_mult_1_multiplication_mult_21_n12,
         my_filter_adder_mult_1_multiplication_mult_21_n11,
         my_filter_adder_mult_1_multiplication_mult_21_n10,
         my_filter_adder_mult_1_multiplication_mult_21_n9,
         my_filter_adder_mult_1_multiplication_mult_21_n8,
         my_filter_adder_mult_1_multiplication_mult_21_n7,
         my_filter_adder_mult_1_multiplication_mult_21_n6,
         my_filter_adder_mult_1_multiplication_mult_21_n5,
         my_filter_adder_mult_1_multiplication_mult_21_n4,
         my_filter_adder_mult_1_multiplication_mult_21_n3,
         my_filter_adder_mult_1_multiplication_mult_21_A2_12_,
         my_filter_adder_mult_1_multiplication_mult_21_A1_0_,
         my_filter_adder_mult_1_multiplication_mult_21_A1_1_,
         my_filter_adder_mult_1_multiplication_mult_21_A1_2_,
         my_filter_adder_mult_1_multiplication_mult_21_A1_3_,
         my_filter_adder_mult_1_multiplication_mult_21_A1_4_,
         my_filter_adder_mult_1_multiplication_mult_21_A1_5_,
         my_filter_adder_mult_1_multiplication_mult_21_A1_6_,
         my_filter_adder_mult_1_multiplication_mult_21_A1_7_,
         my_filter_adder_mult_1_multiplication_mult_21_A1_8_,
         my_filter_adder_mult_1_multiplication_mult_21_A1_9_,
         my_filter_adder_mult_1_multiplication_mult_21_A1_10_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_2__1_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_2__2_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_2__3_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_2__4_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_2__5_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_2__6_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_2__7_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_2__8_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_2__9_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_2__10_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_2__11_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_2__12_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_3__1_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_3__2_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_3__3_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_3__4_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_3__5_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_3__6_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_3__7_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_3__8_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_3__9_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_3__10_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_3__11_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_3__12_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_4__1_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_4__2_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_4__3_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_4__4_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_4__5_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_4__6_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_4__7_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_4__8_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_4__9_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_4__10_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_4__11_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_4__12_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_5__1_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_5__2_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_5__3_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_5__4_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_5__5_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_5__6_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_5__7_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_5__8_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_5__9_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_5__10_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_5__11_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_5__12_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_6__1_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_6__2_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_6__3_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_6__4_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_6__5_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_6__6_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_6__7_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_6__8_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_6__9_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_6__10_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_6__11_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_6__12_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_7__1_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_7__2_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_7__3_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_7__4_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_7__5_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_7__6_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_7__7_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_7__8_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_7__9_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_7__10_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_7__11_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_7__12_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_8__1_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_8__2_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_8__3_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_8__4_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_8__5_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_8__6_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_8__7_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_8__8_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_8__9_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_8__10_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_8__11_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_8__12_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_9__1_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_9__2_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_9__3_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_9__4_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_9__5_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_9__6_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_9__7_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_9__8_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_9__9_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_9__10_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_9__11_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_9__12_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_10__1_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_10__2_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_10__3_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_10__4_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_10__5_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_10__6_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_10__7_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_10__8_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_10__9_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_10__10_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_10__11_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_10__12_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_11__1_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_11__2_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_11__3_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_11__4_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_11__5_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_11__6_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_11__7_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_11__8_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_11__9_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_11__10_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_11__11_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_11__12_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_12__1_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_12__2_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_12__3_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_12__4_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_12__5_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_12__6_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_12__7_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_12__8_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_12__9_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_12__10_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_12__11_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_12__12_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_13__0_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_13__1_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_13__2_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_13__3_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_13__4_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_13__5_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_13__6_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_13__7_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_13__8_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_13__9_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_13__10_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_13__11_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_13__12_,
         my_filter_adder_mult_1_multiplication_mult_21_SUMB_13__13_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_1__0_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_2__0_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_2__1_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_2__2_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_2__3_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_2__4_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_2__5_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_2__6_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_2__7_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_2__8_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_2__9_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_2__10_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_2__11_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_2__12_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_3__0_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_3__1_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_3__2_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_3__3_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_3__4_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_3__5_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_3__6_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_3__7_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_3__8_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_3__9_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_3__10_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_3__11_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_3__12_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_4__0_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_4__1_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_4__2_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_4__3_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_4__4_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_4__5_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_4__6_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_4__7_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_4__8_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_4__9_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_4__10_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_4__11_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_4__12_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_5__0_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_5__1_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_5__2_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_5__3_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_5__4_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_5__5_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_5__6_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_5__7_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_5__8_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_5__9_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_5__10_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_5__11_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_5__12_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_6__0_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_6__1_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_6__2_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_6__3_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_6__4_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_6__5_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_6__6_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_6__7_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_6__8_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_6__9_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_6__10_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_6__11_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_6__12_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_7__0_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_7__1_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_7__2_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_7__3_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_7__4_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_7__5_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_7__6_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_7__7_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_7__8_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_7__9_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_7__10_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_7__11_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_7__12_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_8__0_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_8__1_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_8__2_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_8__3_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_8__4_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_8__5_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_8__6_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_8__7_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_8__8_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_8__9_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_8__10_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_8__11_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_8__12_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_9__0_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_9__1_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_9__2_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_9__3_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_9__4_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_9__5_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_9__6_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_9__7_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_9__8_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_9__9_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_9__10_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_9__11_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_9__12_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_10__0_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_10__1_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_10__2_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_10__3_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_10__4_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_10__5_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_10__6_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_10__7_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_10__8_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_10__9_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_10__10_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_10__11_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_10__12_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_11__0_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_11__1_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_11__2_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_11__3_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_11__4_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_11__5_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_11__6_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_11__7_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_11__8_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_11__9_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_11__10_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_11__11_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_11__12_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_12__0_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_12__1_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_12__2_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_12__3_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_12__4_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_12__5_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_12__6_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_12__7_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_12__8_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_12__9_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_12__10_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_12__11_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_12__12_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_13__0_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_13__1_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_13__2_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_13__3_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_13__4_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_13__5_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_13__6_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_13__7_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_13__8_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_13__9_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_13__10_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_13__11_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_13__12_,
         my_filter_adder_mult_1_multiplication_mult_21_CARRYB_13__13_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_0__2_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_0__3_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_0__4_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_0__5_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_0__6_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_0__7_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_0__8_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_0__9_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_0__10_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_0__11_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_0__12_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_0__13_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_1__1_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_1__2_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_1__3_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_1__4_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_1__5_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_1__6_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_1__7_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_1__8_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_1__9_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_1__10_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_1__11_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_1__12_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_1__13_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_2__0_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_2__1_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_2__2_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_2__3_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_2__4_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_2__5_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_2__6_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_2__7_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_2__8_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_2__9_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_2__10_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_2__11_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_2__12_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_2__13_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_3__0_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_3__1_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_3__2_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_3__3_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_3__4_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_3__5_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_3__6_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_3__7_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_3__8_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_3__9_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_3__10_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_3__11_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_3__12_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_3__13_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_4__0_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_4__1_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_4__2_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_4__3_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_4__4_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_4__5_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_4__6_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_4__7_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_4__8_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_4__9_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_4__10_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_4__11_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_4__12_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_4__13_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_5__0_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_5__1_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_5__2_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_5__3_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_5__4_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_5__5_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_5__6_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_5__7_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_5__8_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_5__9_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_5__10_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_5__11_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_5__12_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_5__13_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_6__0_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_6__1_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_6__2_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_6__3_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_6__4_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_6__5_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_6__6_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_6__7_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_6__8_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_6__9_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_6__10_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_6__11_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_6__12_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_6__13_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_7__0_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_7__1_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_7__2_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_7__3_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_7__4_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_7__5_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_7__6_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_7__7_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_7__8_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_7__9_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_7__10_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_7__11_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_7__12_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_7__13_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_8__0_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_8__1_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_8__2_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_8__3_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_8__4_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_8__5_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_8__6_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_8__7_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_8__8_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_8__9_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_8__10_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_8__11_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_8__12_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_8__13_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_9__0_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_9__1_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_9__2_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_9__3_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_9__4_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_9__5_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_9__6_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_9__7_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_9__8_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_9__9_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_9__10_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_9__11_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_9__12_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_9__13_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_10__0_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_10__1_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_10__2_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_10__3_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_10__4_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_10__5_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_10__6_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_10__7_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_10__8_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_10__9_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_10__10_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_10__11_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_10__12_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_10__13_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_11__0_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_11__1_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_11__2_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_11__3_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_11__4_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_11__5_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_11__6_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_11__7_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_11__8_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_11__9_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_11__10_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_11__11_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_11__12_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_11__13_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_12__0_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_12__1_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_12__2_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_12__3_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_12__4_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_12__5_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_12__6_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_12__7_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_12__8_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_12__9_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_12__10_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_12__11_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_12__12_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_12__13_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_13__0_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_13__1_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_13__2_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_13__3_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_13__4_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_13__5_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_13__6_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_13__7_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_13__8_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_13__9_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_13__10_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_13__11_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_13__12_,
         my_filter_adder_mult_1_multiplication_mult_21_ab_13__13_,
         my_filter_adder_mult_1_multiplication_mult_21_FS_1_n71,
         my_filter_adder_mult_1_multiplication_mult_21_FS_1_n70,
         my_filter_adder_mult_1_multiplication_mult_21_FS_1_n69,
         my_filter_adder_mult_1_multiplication_mult_21_FS_1_n68,
         my_filter_adder_mult_1_multiplication_mult_21_FS_1_n67,
         my_filter_adder_mult_1_multiplication_mult_21_FS_1_n66,
         my_filter_adder_mult_1_multiplication_mult_21_FS_1_n65,
         my_filter_adder_mult_1_multiplication_mult_21_FS_1_n64,
         my_filter_adder_mult_1_multiplication_mult_21_FS_1_n63,
         my_filter_adder_mult_1_multiplication_mult_21_FS_1_n62,
         my_filter_adder_mult_1_multiplication_mult_21_FS_1_n60,
         my_filter_adder_mult_1_multiplication_mult_21_FS_1_n59,
         my_filter_adder_mult_1_multiplication_mult_21_FS_1_n58,
         my_filter_adder_mult_1_multiplication_mult_21_FS_1_n57,
         my_filter_adder_mult_1_multiplication_mult_21_FS_1_n56,
         my_filter_adder_mult_1_multiplication_mult_21_FS_1_n55,
         my_filter_adder_mult_1_multiplication_mult_21_FS_1_n54,
         my_filter_adder_mult_1_multiplication_mult_21_FS_1_n53,
         my_filter_adder_mult_1_multiplication_mult_21_FS_1_n52,
         my_filter_adder_mult_1_multiplication_mult_21_FS_1_n51,
         my_filter_adder_mult_1_multiplication_mult_21_FS_1_n50,
         my_filter_adder_mult_1_multiplication_mult_21_FS_1_n49,
         my_filter_adder_mult_1_multiplication_mult_21_FS_1_n48,
         my_filter_adder_mult_1_multiplication_mult_21_FS_1_n47,
         my_filter_adder_mult_1_multiplication_mult_21_FS_1_n46,
         my_filter_adder_mult_1_multiplication_mult_21_FS_1_n45,
         my_filter_adder_mult_1_multiplication_mult_21_FS_1_n44,
         my_filter_adder_mult_1_multiplication_mult_21_FS_1_n43,
         my_filter_adder_mult_1_multiplication_mult_21_FS_1_n42,
         my_filter_adder_mult_1_multiplication_mult_21_FS_1_n41,
         my_filter_adder_mult_1_multiplication_mult_21_FS_1_n40,
         my_filter_adder_mult_1_multiplication_mult_21_FS_1_n39,
         my_filter_adder_mult_1_multiplication_mult_21_FS_1_n38,
         my_filter_adder_mult_1_multiplication_mult_21_FS_1_n37,
         my_filter_adder_mult_1_multiplication_mult_21_FS_1_n36,
         my_filter_adder_mult_1_multiplication_mult_21_FS_1_n35,
         my_filter_adder_mult_1_multiplication_mult_21_FS_1_n34,
         my_filter_adder_mult_1_multiplication_mult_21_FS_1_n33,
         my_filter_adder_mult_1_multiplication_mult_21_FS_1_n32,
         my_filter_adder_mult_1_multiplication_mult_21_FS_1_n31,
         my_filter_adder_mult_1_multiplication_mult_21_FS_1_n30,
         my_filter_adder_mult_1_multiplication_mult_21_FS_1_n29,
         my_filter_adder_mult_1_multiplication_mult_21_FS_1_n28,
         my_filter_adder_mult_1_multiplication_mult_21_FS_1_n27,
         my_filter_adder_mult_1_multiplication_mult_21_FS_1_n26,
         my_filter_adder_mult_1_multiplication_mult_21_FS_1_n25,
         my_filter_adder_mult_1_multiplication_mult_21_FS_1_n24,
         my_filter_adder_mult_1_multiplication_mult_21_FS_1_n23,
         my_filter_adder_mult_1_multiplication_mult_21_FS_1_n22,
         my_filter_adder_mult_1_multiplication_mult_21_FS_1_n21,
         my_filter_adder_mult_1_multiplication_mult_21_FS_1_n20,
         my_filter_adder_mult_1_multiplication_mult_21_FS_1_n19,
         my_filter_adder_mult_1_multiplication_mult_21_FS_1_n18,
         my_filter_adder_mult_1_multiplication_mult_21_FS_1_n17,
         my_filter_adder_mult_1_multiplication_mult_21_FS_1_n16,
         my_filter_adder_mult_1_multiplication_mult_21_FS_1_n15,
         my_filter_adder_mult_1_multiplication_mult_21_FS_1_n14,
         my_filter_adder_mult_1_multiplication_mult_21_FS_1_n13,
         my_filter_adder_mult_1_addition_add_19_n1,
         my_filter_adder_mult_2_multiplication_mult_21_n113,
         my_filter_adder_mult_2_multiplication_mult_21_n112,
         my_filter_adder_mult_2_multiplication_mult_21_n111,
         my_filter_adder_mult_2_multiplication_mult_21_n110,
         my_filter_adder_mult_2_multiplication_mult_21_n109,
         my_filter_adder_mult_2_multiplication_mult_21_n108,
         my_filter_adder_mult_2_multiplication_mult_21_n107,
         my_filter_adder_mult_2_multiplication_mult_21_n106,
         my_filter_adder_mult_2_multiplication_mult_21_n105,
         my_filter_adder_mult_2_multiplication_mult_21_n104,
         my_filter_adder_mult_2_multiplication_mult_21_n103,
         my_filter_adder_mult_2_multiplication_mult_21_n102,
         my_filter_adder_mult_2_multiplication_mult_21_n101,
         my_filter_adder_mult_2_multiplication_mult_21_n100,
         my_filter_adder_mult_2_multiplication_mult_21_n99,
         my_filter_adder_mult_2_multiplication_mult_21_n98,
         my_filter_adder_mult_2_multiplication_mult_21_n97,
         my_filter_adder_mult_2_multiplication_mult_21_n96,
         my_filter_adder_mult_2_multiplication_mult_21_n95,
         my_filter_adder_mult_2_multiplication_mult_21_n94,
         my_filter_adder_mult_2_multiplication_mult_21_n93,
         my_filter_adder_mult_2_multiplication_mult_21_n92,
         my_filter_adder_mult_2_multiplication_mult_21_n91,
         my_filter_adder_mult_2_multiplication_mult_21_n90,
         my_filter_adder_mult_2_multiplication_mult_21_n89,
         my_filter_adder_mult_2_multiplication_mult_21_n88,
         my_filter_adder_mult_2_multiplication_mult_21_n87,
         my_filter_adder_mult_2_multiplication_mult_21_n86,
         my_filter_adder_mult_2_multiplication_mult_21_n85,
         my_filter_adder_mult_2_multiplication_mult_21_n52,
         my_filter_adder_mult_2_multiplication_mult_21_n51,
         my_filter_adder_mult_2_multiplication_mult_21_n50,
         my_filter_adder_mult_2_multiplication_mult_21_n49,
         my_filter_adder_mult_2_multiplication_mult_21_n48,
         my_filter_adder_mult_2_multiplication_mult_21_n47,
         my_filter_adder_mult_2_multiplication_mult_21_n46,
         my_filter_adder_mult_2_multiplication_mult_21_n45,
         my_filter_adder_mult_2_multiplication_mult_21_n44,
         my_filter_adder_mult_2_multiplication_mult_21_n43,
         my_filter_adder_mult_2_multiplication_mult_21_n42,
         my_filter_adder_mult_2_multiplication_mult_21_n41,
         my_filter_adder_mult_2_multiplication_mult_21_n40,
         my_filter_adder_mult_2_multiplication_mult_21_n39,
         my_filter_adder_mult_2_multiplication_mult_21_n38,
         my_filter_adder_mult_2_multiplication_mult_21_n37,
         my_filter_adder_mult_2_multiplication_mult_21_n36,
         my_filter_adder_mult_2_multiplication_mult_21_n35,
         my_filter_adder_mult_2_multiplication_mult_21_n34,
         my_filter_adder_mult_2_multiplication_mult_21_n33,
         my_filter_adder_mult_2_multiplication_mult_21_n32,
         my_filter_adder_mult_2_multiplication_mult_21_n31,
         my_filter_adder_mult_2_multiplication_mult_21_n30,
         my_filter_adder_mult_2_multiplication_mult_21_n29,
         my_filter_adder_mult_2_multiplication_mult_21_n28,
         my_filter_adder_mult_2_multiplication_mult_21_n27,
         my_filter_adder_mult_2_multiplication_mult_21_n26,
         my_filter_adder_mult_2_multiplication_mult_21_n25,
         my_filter_adder_mult_2_multiplication_mult_21_n24,
         my_filter_adder_mult_2_multiplication_mult_21_n23,
         my_filter_adder_mult_2_multiplication_mult_21_n22,
         my_filter_adder_mult_2_multiplication_mult_21_n21,
         my_filter_adder_mult_2_multiplication_mult_21_n20,
         my_filter_adder_mult_2_multiplication_mult_21_n19,
         my_filter_adder_mult_2_multiplication_mult_21_n18,
         my_filter_adder_mult_2_multiplication_mult_21_n17,
         my_filter_adder_mult_2_multiplication_mult_21_n16,
         my_filter_adder_mult_2_multiplication_mult_21_n15,
         my_filter_adder_mult_2_multiplication_mult_21_n14,
         my_filter_adder_mult_2_multiplication_mult_21_n13,
         my_filter_adder_mult_2_multiplication_mult_21_n12,
         my_filter_adder_mult_2_multiplication_mult_21_n11,
         my_filter_adder_mult_2_multiplication_mult_21_n10,
         my_filter_adder_mult_2_multiplication_mult_21_n9,
         my_filter_adder_mult_2_multiplication_mult_21_n8,
         my_filter_adder_mult_2_multiplication_mult_21_n7,
         my_filter_adder_mult_2_multiplication_mult_21_n6,
         my_filter_adder_mult_2_multiplication_mult_21_n5,
         my_filter_adder_mult_2_multiplication_mult_21_n4,
         my_filter_adder_mult_2_multiplication_mult_21_n3,
         my_filter_adder_mult_2_multiplication_mult_21_A2_12_,
         my_filter_adder_mult_2_multiplication_mult_21_A1_0_,
         my_filter_adder_mult_2_multiplication_mult_21_A1_1_,
         my_filter_adder_mult_2_multiplication_mult_21_A1_2_,
         my_filter_adder_mult_2_multiplication_mult_21_A1_3_,
         my_filter_adder_mult_2_multiplication_mult_21_A1_4_,
         my_filter_adder_mult_2_multiplication_mult_21_A1_5_,
         my_filter_adder_mult_2_multiplication_mult_21_A1_6_,
         my_filter_adder_mult_2_multiplication_mult_21_A1_7_,
         my_filter_adder_mult_2_multiplication_mult_21_A1_8_,
         my_filter_adder_mult_2_multiplication_mult_21_A1_9_,
         my_filter_adder_mult_2_multiplication_mult_21_A1_10_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_2__1_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_2__2_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_2__3_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_2__4_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_2__5_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_2__6_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_2__7_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_2__8_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_2__9_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_2__10_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_2__11_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_2__12_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_3__1_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_3__2_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_3__3_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_3__4_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_3__5_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_3__6_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_3__7_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_3__8_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_3__9_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_3__10_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_3__11_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_3__12_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_4__1_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_4__2_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_4__3_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_4__4_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_4__5_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_4__6_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_4__7_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_4__8_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_4__9_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_4__10_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_4__11_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_4__12_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_5__1_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_5__2_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_5__3_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_5__4_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_5__5_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_5__6_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_5__7_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_5__8_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_5__9_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_5__10_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_5__11_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_5__12_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_6__1_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_6__2_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_6__3_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_6__4_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_6__5_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_6__6_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_6__7_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_6__8_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_6__9_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_6__10_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_6__11_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_6__12_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_7__1_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_7__2_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_7__3_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_7__4_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_7__5_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_7__6_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_7__7_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_7__8_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_7__9_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_7__10_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_7__11_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_7__12_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_8__1_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_8__2_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_8__3_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_8__4_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_8__5_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_8__6_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_8__7_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_8__8_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_8__9_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_8__10_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_8__11_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_8__12_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_9__1_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_9__2_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_9__3_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_9__4_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_9__5_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_9__6_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_9__7_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_9__8_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_9__9_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_9__10_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_9__11_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_9__12_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_10__1_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_10__2_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_10__3_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_10__4_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_10__5_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_10__6_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_10__7_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_10__8_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_10__9_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_10__10_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_10__11_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_10__12_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_11__1_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_11__2_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_11__3_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_11__4_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_11__5_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_11__6_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_11__7_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_11__8_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_11__9_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_11__10_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_11__11_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_11__12_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_12__1_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_12__2_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_12__3_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_12__4_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_12__5_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_12__6_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_12__7_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_12__8_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_12__9_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_12__10_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_12__11_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_12__12_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_13__0_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_13__1_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_13__2_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_13__3_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_13__4_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_13__5_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_13__6_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_13__7_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_13__8_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_13__9_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_13__10_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_13__11_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_13__12_,
         my_filter_adder_mult_2_multiplication_mult_21_SUMB_13__13_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_1__0_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_2__0_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_2__1_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_2__2_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_2__3_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_2__4_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_2__5_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_2__6_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_2__7_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_2__8_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_2__9_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_2__10_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_2__11_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_2__12_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_3__0_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_3__1_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_3__2_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_3__3_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_3__4_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_3__5_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_3__6_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_3__7_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_3__8_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_3__9_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_3__10_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_3__11_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_3__12_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_4__0_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_4__1_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_4__2_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_4__3_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_4__4_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_4__5_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_4__6_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_4__7_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_4__8_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_4__9_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_4__10_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_4__11_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_4__12_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_5__0_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_5__1_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_5__2_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_5__3_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_5__4_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_5__5_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_5__6_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_5__7_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_5__8_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_5__9_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_5__10_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_5__11_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_5__12_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_6__0_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_6__1_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_6__2_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_6__3_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_6__4_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_6__5_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_6__6_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_6__7_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_6__8_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_6__9_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_6__10_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_6__11_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_6__12_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_7__0_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_7__1_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_7__2_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_7__3_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_7__4_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_7__5_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_7__6_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_7__7_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_7__8_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_7__9_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_7__10_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_7__11_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_7__12_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_8__0_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_8__1_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_8__2_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_8__3_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_8__4_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_8__5_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_8__6_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_8__7_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_8__8_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_8__9_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_8__10_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_8__11_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_8__12_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_9__0_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_9__1_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_9__2_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_9__3_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_9__4_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_9__5_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_9__6_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_9__7_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_9__8_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_9__9_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_9__10_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_9__11_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_9__12_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_10__0_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_10__1_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_10__2_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_10__3_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_10__4_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_10__5_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_10__6_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_10__7_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_10__8_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_10__9_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_10__10_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_10__11_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_10__12_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_11__0_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_11__1_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_11__2_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_11__3_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_11__4_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_11__5_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_11__6_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_11__7_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_11__8_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_11__9_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_11__10_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_11__11_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_11__12_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_12__0_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_12__1_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_12__2_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_12__3_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_12__4_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_12__5_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_12__6_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_12__7_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_12__8_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_12__9_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_12__10_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_12__11_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_12__12_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_13__0_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_13__1_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_13__2_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_13__3_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_13__4_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_13__5_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_13__6_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_13__7_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_13__8_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_13__9_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_13__10_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_13__11_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_13__12_,
         my_filter_adder_mult_2_multiplication_mult_21_CARRYB_13__13_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_0__2_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_0__3_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_0__4_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_0__5_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_0__6_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_0__7_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_0__8_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_0__9_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_0__10_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_0__11_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_0__12_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_0__13_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_1__1_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_1__2_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_1__3_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_1__4_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_1__5_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_1__6_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_1__7_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_1__8_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_1__9_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_1__10_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_1__11_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_1__12_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_1__13_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_2__0_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_2__1_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_2__2_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_2__3_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_2__4_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_2__5_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_2__6_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_2__7_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_2__8_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_2__9_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_2__10_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_2__11_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_2__12_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_2__13_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_3__0_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_3__1_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_3__2_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_3__3_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_3__4_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_3__5_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_3__6_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_3__7_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_3__8_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_3__9_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_3__10_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_3__11_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_3__12_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_3__13_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_4__0_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_4__1_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_4__2_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_4__3_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_4__4_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_4__5_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_4__6_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_4__7_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_4__8_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_4__9_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_4__10_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_4__11_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_4__12_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_4__13_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_5__0_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_5__1_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_5__2_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_5__3_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_5__4_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_5__5_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_5__6_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_5__7_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_5__8_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_5__9_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_5__10_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_5__11_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_5__12_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_5__13_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_6__0_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_6__1_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_6__2_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_6__3_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_6__4_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_6__5_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_6__6_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_6__7_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_6__8_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_6__9_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_6__10_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_6__11_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_6__12_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_6__13_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_7__0_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_7__1_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_7__2_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_7__3_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_7__4_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_7__5_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_7__6_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_7__7_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_7__8_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_7__9_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_7__10_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_7__11_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_7__12_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_7__13_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_8__0_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_8__1_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_8__2_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_8__3_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_8__4_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_8__5_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_8__6_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_8__7_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_8__8_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_8__9_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_8__10_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_8__11_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_8__12_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_8__13_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_9__0_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_9__1_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_9__2_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_9__3_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_9__4_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_9__5_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_9__6_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_9__7_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_9__8_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_9__9_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_9__10_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_9__11_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_9__12_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_9__13_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_10__0_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_10__1_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_10__2_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_10__3_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_10__4_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_10__5_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_10__6_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_10__7_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_10__8_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_10__9_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_10__10_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_10__11_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_10__12_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_10__13_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_11__0_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_11__1_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_11__2_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_11__3_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_11__4_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_11__5_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_11__6_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_11__7_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_11__8_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_11__9_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_11__10_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_11__11_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_11__12_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_11__13_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_12__0_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_12__1_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_12__2_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_12__3_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_12__4_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_12__5_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_12__6_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_12__7_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_12__8_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_12__9_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_12__10_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_12__11_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_12__12_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_12__13_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_13__0_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_13__1_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_13__2_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_13__3_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_13__4_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_13__5_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_13__6_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_13__7_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_13__8_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_13__9_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_13__10_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_13__11_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_13__12_,
         my_filter_adder_mult_2_multiplication_mult_21_ab_13__13_,
         my_filter_adder_mult_2_multiplication_mult_21_FS_1_n71,
         my_filter_adder_mult_2_multiplication_mult_21_FS_1_n70,
         my_filter_adder_mult_2_multiplication_mult_21_FS_1_n69,
         my_filter_adder_mult_2_multiplication_mult_21_FS_1_n68,
         my_filter_adder_mult_2_multiplication_mult_21_FS_1_n67,
         my_filter_adder_mult_2_multiplication_mult_21_FS_1_n66,
         my_filter_adder_mult_2_multiplication_mult_21_FS_1_n65,
         my_filter_adder_mult_2_multiplication_mult_21_FS_1_n64,
         my_filter_adder_mult_2_multiplication_mult_21_FS_1_n63,
         my_filter_adder_mult_2_multiplication_mult_21_FS_1_n62,
         my_filter_adder_mult_2_multiplication_mult_21_FS_1_n60,
         my_filter_adder_mult_2_multiplication_mult_21_FS_1_n59,
         my_filter_adder_mult_2_multiplication_mult_21_FS_1_n58,
         my_filter_adder_mult_2_multiplication_mult_21_FS_1_n57,
         my_filter_adder_mult_2_multiplication_mult_21_FS_1_n56,
         my_filter_adder_mult_2_multiplication_mult_21_FS_1_n55,
         my_filter_adder_mult_2_multiplication_mult_21_FS_1_n54,
         my_filter_adder_mult_2_multiplication_mult_21_FS_1_n53,
         my_filter_adder_mult_2_multiplication_mult_21_FS_1_n52,
         my_filter_adder_mult_2_multiplication_mult_21_FS_1_n51,
         my_filter_adder_mult_2_multiplication_mult_21_FS_1_n50,
         my_filter_adder_mult_2_multiplication_mult_21_FS_1_n49,
         my_filter_adder_mult_2_multiplication_mult_21_FS_1_n48,
         my_filter_adder_mult_2_multiplication_mult_21_FS_1_n47,
         my_filter_adder_mult_2_multiplication_mult_21_FS_1_n46,
         my_filter_adder_mult_2_multiplication_mult_21_FS_1_n45,
         my_filter_adder_mult_2_multiplication_mult_21_FS_1_n44,
         my_filter_adder_mult_2_multiplication_mult_21_FS_1_n43,
         my_filter_adder_mult_2_multiplication_mult_21_FS_1_n42,
         my_filter_adder_mult_2_multiplication_mult_21_FS_1_n41,
         my_filter_adder_mult_2_multiplication_mult_21_FS_1_n40,
         my_filter_adder_mult_2_multiplication_mult_21_FS_1_n39,
         my_filter_adder_mult_2_multiplication_mult_21_FS_1_n38,
         my_filter_adder_mult_2_multiplication_mult_21_FS_1_n37,
         my_filter_adder_mult_2_multiplication_mult_21_FS_1_n36,
         my_filter_adder_mult_2_multiplication_mult_21_FS_1_n35,
         my_filter_adder_mult_2_multiplication_mult_21_FS_1_n34,
         my_filter_adder_mult_2_multiplication_mult_21_FS_1_n33,
         my_filter_adder_mult_2_multiplication_mult_21_FS_1_n32,
         my_filter_adder_mult_2_multiplication_mult_21_FS_1_n31,
         my_filter_adder_mult_2_multiplication_mult_21_FS_1_n30,
         my_filter_adder_mult_2_multiplication_mult_21_FS_1_n29,
         my_filter_adder_mult_2_multiplication_mult_21_FS_1_n28,
         my_filter_adder_mult_2_multiplication_mult_21_FS_1_n27,
         my_filter_adder_mult_2_multiplication_mult_21_FS_1_n26,
         my_filter_adder_mult_2_multiplication_mult_21_FS_1_n25,
         my_filter_adder_mult_2_multiplication_mult_21_FS_1_n24,
         my_filter_adder_mult_2_multiplication_mult_21_FS_1_n23,
         my_filter_adder_mult_2_multiplication_mult_21_FS_1_n22,
         my_filter_adder_mult_2_multiplication_mult_21_FS_1_n21,
         my_filter_adder_mult_2_multiplication_mult_21_FS_1_n20,
         my_filter_adder_mult_2_multiplication_mult_21_FS_1_n19,
         my_filter_adder_mult_2_multiplication_mult_21_FS_1_n18,
         my_filter_adder_mult_2_multiplication_mult_21_FS_1_n17,
         my_filter_adder_mult_2_multiplication_mult_21_FS_1_n16,
         my_filter_adder_mult_2_multiplication_mult_21_FS_1_n15,
         my_filter_adder_mult_2_multiplication_mult_21_FS_1_n14,
         my_filter_adder_mult_2_multiplication_mult_21_FS_1_n13,
         my_filter_adder_mult_2_addition_add_19_n1,
         my_filter_adder_mult_3_multiplication_mult_21_n113,
         my_filter_adder_mult_3_multiplication_mult_21_n112,
         my_filter_adder_mult_3_multiplication_mult_21_n111,
         my_filter_adder_mult_3_multiplication_mult_21_n110,
         my_filter_adder_mult_3_multiplication_mult_21_n109,
         my_filter_adder_mult_3_multiplication_mult_21_n108,
         my_filter_adder_mult_3_multiplication_mult_21_n107,
         my_filter_adder_mult_3_multiplication_mult_21_n106,
         my_filter_adder_mult_3_multiplication_mult_21_n105,
         my_filter_adder_mult_3_multiplication_mult_21_n104,
         my_filter_adder_mult_3_multiplication_mult_21_n103,
         my_filter_adder_mult_3_multiplication_mult_21_n102,
         my_filter_adder_mult_3_multiplication_mult_21_n101,
         my_filter_adder_mult_3_multiplication_mult_21_n100,
         my_filter_adder_mult_3_multiplication_mult_21_n99,
         my_filter_adder_mult_3_multiplication_mult_21_n98,
         my_filter_adder_mult_3_multiplication_mult_21_n97,
         my_filter_adder_mult_3_multiplication_mult_21_n96,
         my_filter_adder_mult_3_multiplication_mult_21_n95,
         my_filter_adder_mult_3_multiplication_mult_21_n94,
         my_filter_adder_mult_3_multiplication_mult_21_n93,
         my_filter_adder_mult_3_multiplication_mult_21_n92,
         my_filter_adder_mult_3_multiplication_mult_21_n91,
         my_filter_adder_mult_3_multiplication_mult_21_n90,
         my_filter_adder_mult_3_multiplication_mult_21_n89,
         my_filter_adder_mult_3_multiplication_mult_21_n88,
         my_filter_adder_mult_3_multiplication_mult_21_n87,
         my_filter_adder_mult_3_multiplication_mult_21_n86,
         my_filter_adder_mult_3_multiplication_mult_21_n85,
         my_filter_adder_mult_3_multiplication_mult_21_n52,
         my_filter_adder_mult_3_multiplication_mult_21_n51,
         my_filter_adder_mult_3_multiplication_mult_21_n50,
         my_filter_adder_mult_3_multiplication_mult_21_n49,
         my_filter_adder_mult_3_multiplication_mult_21_n48,
         my_filter_adder_mult_3_multiplication_mult_21_n47,
         my_filter_adder_mult_3_multiplication_mult_21_n46,
         my_filter_adder_mult_3_multiplication_mult_21_n45,
         my_filter_adder_mult_3_multiplication_mult_21_n44,
         my_filter_adder_mult_3_multiplication_mult_21_n43,
         my_filter_adder_mult_3_multiplication_mult_21_n42,
         my_filter_adder_mult_3_multiplication_mult_21_n41,
         my_filter_adder_mult_3_multiplication_mult_21_n40,
         my_filter_adder_mult_3_multiplication_mult_21_n39,
         my_filter_adder_mult_3_multiplication_mult_21_n38,
         my_filter_adder_mult_3_multiplication_mult_21_n37,
         my_filter_adder_mult_3_multiplication_mult_21_n36,
         my_filter_adder_mult_3_multiplication_mult_21_n35,
         my_filter_adder_mult_3_multiplication_mult_21_n34,
         my_filter_adder_mult_3_multiplication_mult_21_n33,
         my_filter_adder_mult_3_multiplication_mult_21_n32,
         my_filter_adder_mult_3_multiplication_mult_21_n31,
         my_filter_adder_mult_3_multiplication_mult_21_n30,
         my_filter_adder_mult_3_multiplication_mult_21_n29,
         my_filter_adder_mult_3_multiplication_mult_21_n28,
         my_filter_adder_mult_3_multiplication_mult_21_n27,
         my_filter_adder_mult_3_multiplication_mult_21_n26,
         my_filter_adder_mult_3_multiplication_mult_21_n25,
         my_filter_adder_mult_3_multiplication_mult_21_n24,
         my_filter_adder_mult_3_multiplication_mult_21_n23,
         my_filter_adder_mult_3_multiplication_mult_21_n22,
         my_filter_adder_mult_3_multiplication_mult_21_n21,
         my_filter_adder_mult_3_multiplication_mult_21_n20,
         my_filter_adder_mult_3_multiplication_mult_21_n19,
         my_filter_adder_mult_3_multiplication_mult_21_n18,
         my_filter_adder_mult_3_multiplication_mult_21_n17,
         my_filter_adder_mult_3_multiplication_mult_21_n16,
         my_filter_adder_mult_3_multiplication_mult_21_n15,
         my_filter_adder_mult_3_multiplication_mult_21_n14,
         my_filter_adder_mult_3_multiplication_mult_21_n13,
         my_filter_adder_mult_3_multiplication_mult_21_n12,
         my_filter_adder_mult_3_multiplication_mult_21_n11,
         my_filter_adder_mult_3_multiplication_mult_21_n10,
         my_filter_adder_mult_3_multiplication_mult_21_n9,
         my_filter_adder_mult_3_multiplication_mult_21_n8,
         my_filter_adder_mult_3_multiplication_mult_21_n7,
         my_filter_adder_mult_3_multiplication_mult_21_n6,
         my_filter_adder_mult_3_multiplication_mult_21_n5,
         my_filter_adder_mult_3_multiplication_mult_21_n4,
         my_filter_adder_mult_3_multiplication_mult_21_n3,
         my_filter_adder_mult_3_multiplication_mult_21_A2_12_,
         my_filter_adder_mult_3_multiplication_mult_21_A1_0_,
         my_filter_adder_mult_3_multiplication_mult_21_A1_1_,
         my_filter_adder_mult_3_multiplication_mult_21_A1_2_,
         my_filter_adder_mult_3_multiplication_mult_21_A1_3_,
         my_filter_adder_mult_3_multiplication_mult_21_A1_4_,
         my_filter_adder_mult_3_multiplication_mult_21_A1_5_,
         my_filter_adder_mult_3_multiplication_mult_21_A1_6_,
         my_filter_adder_mult_3_multiplication_mult_21_A1_7_,
         my_filter_adder_mult_3_multiplication_mult_21_A1_8_,
         my_filter_adder_mult_3_multiplication_mult_21_A1_9_,
         my_filter_adder_mult_3_multiplication_mult_21_A1_10_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_2__1_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_2__2_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_2__3_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_2__4_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_2__5_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_2__6_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_2__7_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_2__8_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_2__9_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_2__10_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_2__11_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_2__12_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_3__1_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_3__2_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_3__3_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_3__4_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_3__5_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_3__6_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_3__7_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_3__8_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_3__9_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_3__10_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_3__11_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_3__12_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_4__1_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_4__2_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_4__3_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_4__4_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_4__5_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_4__6_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_4__7_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_4__8_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_4__9_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_4__10_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_4__11_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_4__12_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_5__1_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_5__2_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_5__3_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_5__4_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_5__5_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_5__6_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_5__7_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_5__8_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_5__9_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_5__10_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_5__11_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_5__12_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_6__1_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_6__2_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_6__3_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_6__4_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_6__5_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_6__6_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_6__7_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_6__8_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_6__9_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_6__10_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_6__11_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_6__12_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_7__1_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_7__2_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_7__3_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_7__4_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_7__5_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_7__6_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_7__7_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_7__8_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_7__9_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_7__10_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_7__11_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_7__12_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_8__1_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_8__2_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_8__3_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_8__4_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_8__5_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_8__6_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_8__7_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_8__8_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_8__9_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_8__10_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_8__11_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_8__12_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_9__1_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_9__2_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_9__3_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_9__4_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_9__5_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_9__6_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_9__7_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_9__8_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_9__9_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_9__10_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_9__11_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_9__12_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_10__1_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_10__2_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_10__3_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_10__4_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_10__5_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_10__6_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_10__7_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_10__8_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_10__9_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_10__10_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_10__11_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_10__12_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_11__1_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_11__2_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_11__3_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_11__4_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_11__5_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_11__6_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_11__7_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_11__8_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_11__9_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_11__10_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_11__11_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_11__12_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_12__1_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_12__2_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_12__3_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_12__4_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_12__5_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_12__6_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_12__7_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_12__8_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_12__9_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_12__10_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_12__11_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_12__12_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_13__0_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_13__1_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_13__2_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_13__3_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_13__4_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_13__5_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_13__6_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_13__7_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_13__8_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_13__9_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_13__10_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_13__11_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_13__12_,
         my_filter_adder_mult_3_multiplication_mult_21_SUMB_13__13_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_1__0_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_2__0_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_2__1_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_2__2_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_2__3_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_2__4_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_2__5_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_2__6_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_2__7_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_2__8_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_2__9_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_2__10_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_2__11_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_2__12_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_3__0_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_3__1_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_3__2_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_3__3_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_3__4_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_3__5_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_3__6_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_3__7_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_3__8_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_3__9_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_3__10_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_3__11_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_3__12_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_4__0_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_4__1_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_4__2_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_4__3_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_4__4_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_4__5_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_4__6_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_4__7_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_4__8_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_4__9_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_4__10_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_4__11_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_4__12_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_5__0_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_5__1_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_5__2_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_5__3_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_5__4_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_5__5_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_5__6_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_5__7_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_5__8_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_5__9_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_5__10_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_5__11_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_5__12_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_6__0_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_6__1_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_6__2_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_6__3_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_6__4_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_6__5_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_6__6_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_6__7_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_6__8_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_6__9_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_6__10_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_6__11_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_6__12_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_7__0_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_7__1_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_7__2_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_7__3_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_7__4_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_7__5_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_7__6_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_7__7_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_7__8_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_7__9_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_7__10_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_7__11_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_7__12_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_8__0_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_8__1_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_8__2_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_8__3_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_8__4_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_8__5_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_8__6_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_8__7_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_8__8_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_8__9_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_8__10_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_8__11_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_8__12_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_9__0_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_9__1_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_9__2_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_9__3_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_9__4_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_9__5_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_9__6_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_9__7_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_9__8_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_9__9_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_9__10_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_9__11_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_9__12_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_10__0_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_10__1_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_10__2_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_10__3_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_10__4_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_10__5_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_10__6_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_10__7_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_10__8_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_10__9_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_10__10_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_10__11_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_10__12_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_11__0_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_11__1_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_11__2_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_11__3_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_11__4_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_11__5_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_11__6_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_11__7_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_11__8_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_11__9_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_11__10_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_11__11_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_11__12_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_12__0_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_12__1_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_12__2_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_12__3_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_12__4_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_12__5_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_12__6_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_12__7_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_12__8_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_12__9_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_12__10_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_12__11_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_12__12_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_13__0_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_13__1_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_13__2_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_13__3_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_13__4_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_13__5_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_13__6_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_13__7_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_13__8_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_13__9_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_13__10_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_13__11_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_13__12_,
         my_filter_adder_mult_3_multiplication_mult_21_CARRYB_13__13_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_0__2_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_0__3_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_0__4_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_0__5_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_0__6_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_0__7_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_0__8_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_0__9_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_0__10_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_0__11_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_0__12_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_0__13_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_1__1_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_1__2_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_1__3_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_1__4_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_1__5_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_1__6_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_1__7_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_1__8_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_1__9_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_1__10_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_1__11_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_1__12_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_1__13_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_2__0_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_2__1_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_2__2_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_2__3_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_2__4_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_2__5_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_2__6_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_2__7_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_2__8_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_2__9_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_2__10_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_2__11_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_2__12_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_2__13_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_3__0_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_3__1_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_3__2_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_3__3_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_3__4_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_3__5_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_3__6_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_3__7_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_3__8_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_3__9_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_3__10_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_3__11_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_3__12_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_3__13_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_4__0_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_4__1_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_4__2_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_4__3_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_4__4_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_4__5_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_4__6_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_4__7_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_4__8_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_4__9_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_4__10_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_4__11_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_4__12_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_4__13_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_5__0_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_5__1_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_5__2_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_5__3_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_5__4_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_5__5_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_5__6_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_5__7_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_5__8_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_5__9_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_5__10_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_5__11_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_5__12_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_5__13_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_6__0_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_6__1_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_6__2_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_6__3_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_6__4_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_6__5_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_6__6_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_6__7_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_6__8_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_6__9_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_6__10_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_6__11_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_6__12_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_6__13_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_7__0_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_7__1_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_7__2_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_7__3_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_7__4_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_7__5_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_7__6_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_7__7_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_7__8_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_7__9_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_7__10_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_7__11_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_7__12_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_7__13_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_8__0_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_8__1_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_8__2_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_8__3_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_8__4_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_8__5_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_8__6_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_8__7_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_8__8_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_8__9_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_8__10_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_8__11_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_8__12_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_8__13_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_9__0_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_9__1_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_9__2_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_9__3_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_9__4_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_9__5_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_9__6_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_9__7_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_9__8_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_9__9_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_9__10_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_9__11_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_9__12_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_9__13_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_10__0_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_10__1_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_10__2_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_10__3_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_10__4_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_10__5_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_10__6_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_10__7_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_10__8_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_10__9_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_10__10_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_10__11_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_10__12_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_10__13_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_11__0_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_11__1_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_11__2_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_11__3_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_11__4_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_11__5_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_11__6_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_11__7_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_11__8_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_11__9_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_11__10_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_11__11_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_11__12_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_11__13_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_12__0_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_12__1_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_12__2_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_12__3_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_12__4_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_12__5_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_12__6_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_12__7_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_12__8_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_12__9_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_12__10_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_12__11_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_12__12_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_12__13_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_13__0_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_13__1_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_13__2_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_13__3_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_13__4_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_13__5_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_13__6_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_13__7_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_13__8_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_13__9_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_13__10_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_13__11_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_13__12_,
         my_filter_adder_mult_3_multiplication_mult_21_ab_13__13_,
         my_filter_adder_mult_3_multiplication_mult_21_FS_1_n71,
         my_filter_adder_mult_3_multiplication_mult_21_FS_1_n70,
         my_filter_adder_mult_3_multiplication_mult_21_FS_1_n69,
         my_filter_adder_mult_3_multiplication_mult_21_FS_1_n68,
         my_filter_adder_mult_3_multiplication_mult_21_FS_1_n67,
         my_filter_adder_mult_3_multiplication_mult_21_FS_1_n66,
         my_filter_adder_mult_3_multiplication_mult_21_FS_1_n65,
         my_filter_adder_mult_3_multiplication_mult_21_FS_1_n64,
         my_filter_adder_mult_3_multiplication_mult_21_FS_1_n63,
         my_filter_adder_mult_3_multiplication_mult_21_FS_1_n62,
         my_filter_adder_mult_3_multiplication_mult_21_FS_1_n60,
         my_filter_adder_mult_3_multiplication_mult_21_FS_1_n59,
         my_filter_adder_mult_3_multiplication_mult_21_FS_1_n58,
         my_filter_adder_mult_3_multiplication_mult_21_FS_1_n57,
         my_filter_adder_mult_3_multiplication_mult_21_FS_1_n56,
         my_filter_adder_mult_3_multiplication_mult_21_FS_1_n55,
         my_filter_adder_mult_3_multiplication_mult_21_FS_1_n54,
         my_filter_adder_mult_3_multiplication_mult_21_FS_1_n53,
         my_filter_adder_mult_3_multiplication_mult_21_FS_1_n52,
         my_filter_adder_mult_3_multiplication_mult_21_FS_1_n51,
         my_filter_adder_mult_3_multiplication_mult_21_FS_1_n50,
         my_filter_adder_mult_3_multiplication_mult_21_FS_1_n49,
         my_filter_adder_mult_3_multiplication_mult_21_FS_1_n48,
         my_filter_adder_mult_3_multiplication_mult_21_FS_1_n47,
         my_filter_adder_mult_3_multiplication_mult_21_FS_1_n46,
         my_filter_adder_mult_3_multiplication_mult_21_FS_1_n45,
         my_filter_adder_mult_3_multiplication_mult_21_FS_1_n44,
         my_filter_adder_mult_3_multiplication_mult_21_FS_1_n43,
         my_filter_adder_mult_3_multiplication_mult_21_FS_1_n42,
         my_filter_adder_mult_3_multiplication_mult_21_FS_1_n41,
         my_filter_adder_mult_3_multiplication_mult_21_FS_1_n40,
         my_filter_adder_mult_3_multiplication_mult_21_FS_1_n39,
         my_filter_adder_mult_3_multiplication_mult_21_FS_1_n38,
         my_filter_adder_mult_3_multiplication_mult_21_FS_1_n37,
         my_filter_adder_mult_3_multiplication_mult_21_FS_1_n36,
         my_filter_adder_mult_3_multiplication_mult_21_FS_1_n35,
         my_filter_adder_mult_3_multiplication_mult_21_FS_1_n34,
         my_filter_adder_mult_3_multiplication_mult_21_FS_1_n33,
         my_filter_adder_mult_3_multiplication_mult_21_FS_1_n32,
         my_filter_adder_mult_3_multiplication_mult_21_FS_1_n31,
         my_filter_adder_mult_3_multiplication_mult_21_FS_1_n30,
         my_filter_adder_mult_3_multiplication_mult_21_FS_1_n29,
         my_filter_adder_mult_3_multiplication_mult_21_FS_1_n28,
         my_filter_adder_mult_3_multiplication_mult_21_FS_1_n27,
         my_filter_adder_mult_3_multiplication_mult_21_FS_1_n26,
         my_filter_adder_mult_3_multiplication_mult_21_FS_1_n25,
         my_filter_adder_mult_3_multiplication_mult_21_FS_1_n24,
         my_filter_adder_mult_3_multiplication_mult_21_FS_1_n23,
         my_filter_adder_mult_3_multiplication_mult_21_FS_1_n22,
         my_filter_adder_mult_3_multiplication_mult_21_FS_1_n21,
         my_filter_adder_mult_3_multiplication_mult_21_FS_1_n20,
         my_filter_adder_mult_3_multiplication_mult_21_FS_1_n19,
         my_filter_adder_mult_3_multiplication_mult_21_FS_1_n18,
         my_filter_adder_mult_3_multiplication_mult_21_FS_1_n17,
         my_filter_adder_mult_3_multiplication_mult_21_FS_1_n16,
         my_filter_adder_mult_3_multiplication_mult_21_FS_1_n15,
         my_filter_adder_mult_3_multiplication_mult_21_FS_1_n14,
         my_filter_adder_mult_3_multiplication_mult_21_FS_1_n13,
         my_filter_adder_mult_3_addition_add_19_n1,
         my_filter_adder_mult_4_multiplication_mult_21_n113,
         my_filter_adder_mult_4_multiplication_mult_21_n112,
         my_filter_adder_mult_4_multiplication_mult_21_n111,
         my_filter_adder_mult_4_multiplication_mult_21_n110,
         my_filter_adder_mult_4_multiplication_mult_21_n109,
         my_filter_adder_mult_4_multiplication_mult_21_n108,
         my_filter_adder_mult_4_multiplication_mult_21_n107,
         my_filter_adder_mult_4_multiplication_mult_21_n106,
         my_filter_adder_mult_4_multiplication_mult_21_n105,
         my_filter_adder_mult_4_multiplication_mult_21_n104,
         my_filter_adder_mult_4_multiplication_mult_21_n103,
         my_filter_adder_mult_4_multiplication_mult_21_n102,
         my_filter_adder_mult_4_multiplication_mult_21_n101,
         my_filter_adder_mult_4_multiplication_mult_21_n100,
         my_filter_adder_mult_4_multiplication_mult_21_n99,
         my_filter_adder_mult_4_multiplication_mult_21_n98,
         my_filter_adder_mult_4_multiplication_mult_21_n97,
         my_filter_adder_mult_4_multiplication_mult_21_n96,
         my_filter_adder_mult_4_multiplication_mult_21_n95,
         my_filter_adder_mult_4_multiplication_mult_21_n94,
         my_filter_adder_mult_4_multiplication_mult_21_n93,
         my_filter_adder_mult_4_multiplication_mult_21_n92,
         my_filter_adder_mult_4_multiplication_mult_21_n91,
         my_filter_adder_mult_4_multiplication_mult_21_n90,
         my_filter_adder_mult_4_multiplication_mult_21_n89,
         my_filter_adder_mult_4_multiplication_mult_21_n88,
         my_filter_adder_mult_4_multiplication_mult_21_n87,
         my_filter_adder_mult_4_multiplication_mult_21_n86,
         my_filter_adder_mult_4_multiplication_mult_21_n85,
         my_filter_adder_mult_4_multiplication_mult_21_n52,
         my_filter_adder_mult_4_multiplication_mult_21_n51,
         my_filter_adder_mult_4_multiplication_mult_21_n50,
         my_filter_adder_mult_4_multiplication_mult_21_n49,
         my_filter_adder_mult_4_multiplication_mult_21_n48,
         my_filter_adder_mult_4_multiplication_mult_21_n47,
         my_filter_adder_mult_4_multiplication_mult_21_n46,
         my_filter_adder_mult_4_multiplication_mult_21_n45,
         my_filter_adder_mult_4_multiplication_mult_21_n44,
         my_filter_adder_mult_4_multiplication_mult_21_n43,
         my_filter_adder_mult_4_multiplication_mult_21_n42,
         my_filter_adder_mult_4_multiplication_mult_21_n41,
         my_filter_adder_mult_4_multiplication_mult_21_n40,
         my_filter_adder_mult_4_multiplication_mult_21_n39,
         my_filter_adder_mult_4_multiplication_mult_21_n38,
         my_filter_adder_mult_4_multiplication_mult_21_n37,
         my_filter_adder_mult_4_multiplication_mult_21_n36,
         my_filter_adder_mult_4_multiplication_mult_21_n35,
         my_filter_adder_mult_4_multiplication_mult_21_n34,
         my_filter_adder_mult_4_multiplication_mult_21_n33,
         my_filter_adder_mult_4_multiplication_mult_21_n32,
         my_filter_adder_mult_4_multiplication_mult_21_n31,
         my_filter_adder_mult_4_multiplication_mult_21_n30,
         my_filter_adder_mult_4_multiplication_mult_21_n29,
         my_filter_adder_mult_4_multiplication_mult_21_n28,
         my_filter_adder_mult_4_multiplication_mult_21_n27,
         my_filter_adder_mult_4_multiplication_mult_21_n26,
         my_filter_adder_mult_4_multiplication_mult_21_n25,
         my_filter_adder_mult_4_multiplication_mult_21_n24,
         my_filter_adder_mult_4_multiplication_mult_21_n23,
         my_filter_adder_mult_4_multiplication_mult_21_n22,
         my_filter_adder_mult_4_multiplication_mult_21_n21,
         my_filter_adder_mult_4_multiplication_mult_21_n20,
         my_filter_adder_mult_4_multiplication_mult_21_n19,
         my_filter_adder_mult_4_multiplication_mult_21_n18,
         my_filter_adder_mult_4_multiplication_mult_21_n17,
         my_filter_adder_mult_4_multiplication_mult_21_n16,
         my_filter_adder_mult_4_multiplication_mult_21_n15,
         my_filter_adder_mult_4_multiplication_mult_21_n14,
         my_filter_adder_mult_4_multiplication_mult_21_n13,
         my_filter_adder_mult_4_multiplication_mult_21_n12,
         my_filter_adder_mult_4_multiplication_mult_21_n11,
         my_filter_adder_mult_4_multiplication_mult_21_n10,
         my_filter_adder_mult_4_multiplication_mult_21_n9,
         my_filter_adder_mult_4_multiplication_mult_21_n8,
         my_filter_adder_mult_4_multiplication_mult_21_n7,
         my_filter_adder_mult_4_multiplication_mult_21_n6,
         my_filter_adder_mult_4_multiplication_mult_21_n5,
         my_filter_adder_mult_4_multiplication_mult_21_n4,
         my_filter_adder_mult_4_multiplication_mult_21_n3,
         my_filter_adder_mult_4_multiplication_mult_21_A2_12_,
         my_filter_adder_mult_4_multiplication_mult_21_A1_0_,
         my_filter_adder_mult_4_multiplication_mult_21_A1_1_,
         my_filter_adder_mult_4_multiplication_mult_21_A1_2_,
         my_filter_adder_mult_4_multiplication_mult_21_A1_3_,
         my_filter_adder_mult_4_multiplication_mult_21_A1_4_,
         my_filter_adder_mult_4_multiplication_mult_21_A1_5_,
         my_filter_adder_mult_4_multiplication_mult_21_A1_6_,
         my_filter_adder_mult_4_multiplication_mult_21_A1_7_,
         my_filter_adder_mult_4_multiplication_mult_21_A1_8_,
         my_filter_adder_mult_4_multiplication_mult_21_A1_9_,
         my_filter_adder_mult_4_multiplication_mult_21_A1_10_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_2__1_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_2__2_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_2__3_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_2__4_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_2__5_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_2__6_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_2__7_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_2__8_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_2__9_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_2__10_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_2__11_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_2__12_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_3__1_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_3__2_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_3__3_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_3__4_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_3__5_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_3__6_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_3__7_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_3__8_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_3__9_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_3__10_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_3__11_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_3__12_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_4__1_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_4__2_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_4__3_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_4__4_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_4__5_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_4__6_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_4__7_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_4__8_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_4__9_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_4__10_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_4__11_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_4__12_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_5__1_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_5__2_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_5__3_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_5__4_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_5__5_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_5__6_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_5__7_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_5__8_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_5__9_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_5__10_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_5__11_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_5__12_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_6__1_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_6__2_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_6__3_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_6__4_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_6__5_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_6__6_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_6__7_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_6__8_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_6__9_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_6__10_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_6__11_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_6__12_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_7__1_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_7__2_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_7__3_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_7__4_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_7__5_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_7__6_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_7__7_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_7__8_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_7__9_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_7__10_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_7__11_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_7__12_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_8__1_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_8__2_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_8__3_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_8__4_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_8__5_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_8__6_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_8__7_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_8__8_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_8__9_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_8__10_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_8__11_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_8__12_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_9__1_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_9__2_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_9__3_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_9__4_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_9__5_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_9__6_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_9__7_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_9__8_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_9__9_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_9__10_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_9__11_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_9__12_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_10__1_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_10__2_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_10__3_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_10__4_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_10__5_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_10__6_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_10__7_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_10__8_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_10__9_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_10__10_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_10__11_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_10__12_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_11__1_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_11__2_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_11__3_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_11__4_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_11__5_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_11__6_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_11__7_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_11__8_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_11__9_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_11__10_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_11__11_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_11__12_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_12__1_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_12__2_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_12__3_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_12__4_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_12__5_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_12__6_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_12__7_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_12__8_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_12__9_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_12__10_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_12__11_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_12__12_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_13__0_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_13__1_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_13__2_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_13__3_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_13__4_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_13__5_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_13__6_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_13__7_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_13__8_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_13__9_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_13__10_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_13__11_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_13__12_,
         my_filter_adder_mult_4_multiplication_mult_21_SUMB_13__13_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_1__0_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_2__0_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_2__1_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_2__2_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_2__3_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_2__4_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_2__5_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_2__6_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_2__7_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_2__8_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_2__9_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_2__10_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_2__11_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_2__12_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_3__0_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_3__1_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_3__2_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_3__3_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_3__4_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_3__5_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_3__6_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_3__7_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_3__8_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_3__9_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_3__10_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_3__11_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_3__12_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_4__0_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_4__1_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_4__2_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_4__3_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_4__4_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_4__5_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_4__6_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_4__7_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_4__8_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_4__9_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_4__10_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_4__11_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_4__12_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_5__0_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_5__1_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_5__2_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_5__3_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_5__4_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_5__5_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_5__6_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_5__7_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_5__8_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_5__9_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_5__10_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_5__11_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_5__12_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_6__0_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_6__1_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_6__2_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_6__3_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_6__4_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_6__5_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_6__6_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_6__7_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_6__8_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_6__9_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_6__10_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_6__11_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_6__12_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_7__0_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_7__1_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_7__2_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_7__3_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_7__4_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_7__5_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_7__6_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_7__7_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_7__8_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_7__9_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_7__10_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_7__11_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_7__12_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_8__0_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_8__1_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_8__2_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_8__3_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_8__4_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_8__5_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_8__6_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_8__7_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_8__8_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_8__9_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_8__10_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_8__11_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_8__12_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_9__0_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_9__1_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_9__2_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_9__3_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_9__4_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_9__5_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_9__6_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_9__7_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_9__8_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_9__9_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_9__10_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_9__11_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_9__12_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_10__0_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_10__1_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_10__2_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_10__3_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_10__4_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_10__5_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_10__6_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_10__7_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_10__8_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_10__9_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_10__10_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_10__11_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_10__12_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_11__0_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_11__1_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_11__2_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_11__3_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_11__4_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_11__5_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_11__6_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_11__7_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_11__8_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_11__9_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_11__10_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_11__11_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_11__12_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_12__0_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_12__1_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_12__2_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_12__3_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_12__4_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_12__5_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_12__6_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_12__7_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_12__8_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_12__9_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_12__10_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_12__11_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_12__12_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_13__0_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_13__1_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_13__2_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_13__3_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_13__4_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_13__5_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_13__6_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_13__7_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_13__8_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_13__9_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_13__10_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_13__11_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_13__12_,
         my_filter_adder_mult_4_multiplication_mult_21_CARRYB_13__13_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_0__2_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_0__3_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_0__4_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_0__5_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_0__6_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_0__7_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_0__8_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_0__9_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_0__10_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_0__11_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_0__12_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_0__13_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_1__1_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_1__2_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_1__3_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_1__4_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_1__5_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_1__6_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_1__7_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_1__8_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_1__9_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_1__10_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_1__11_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_1__12_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_1__13_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_2__0_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_2__1_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_2__2_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_2__3_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_2__4_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_2__5_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_2__6_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_2__7_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_2__8_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_2__9_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_2__10_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_2__11_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_2__12_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_2__13_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_3__0_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_3__1_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_3__2_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_3__3_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_3__4_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_3__5_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_3__6_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_3__7_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_3__8_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_3__9_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_3__10_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_3__11_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_3__12_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_3__13_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_4__0_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_4__1_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_4__2_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_4__3_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_4__4_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_4__5_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_4__6_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_4__7_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_4__8_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_4__9_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_4__10_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_4__11_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_4__12_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_4__13_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_5__0_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_5__1_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_5__2_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_5__3_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_5__4_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_5__5_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_5__6_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_5__7_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_5__8_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_5__9_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_5__10_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_5__11_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_5__12_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_5__13_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_6__0_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_6__1_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_6__2_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_6__3_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_6__4_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_6__5_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_6__6_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_6__7_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_6__8_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_6__9_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_6__10_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_6__11_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_6__12_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_6__13_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_7__0_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_7__1_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_7__2_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_7__3_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_7__4_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_7__5_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_7__6_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_7__7_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_7__8_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_7__9_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_7__10_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_7__11_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_7__12_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_7__13_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_8__0_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_8__1_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_8__2_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_8__3_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_8__4_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_8__5_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_8__6_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_8__7_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_8__8_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_8__9_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_8__10_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_8__11_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_8__12_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_8__13_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_9__0_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_9__1_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_9__2_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_9__3_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_9__4_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_9__5_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_9__6_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_9__7_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_9__8_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_9__9_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_9__10_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_9__11_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_9__12_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_9__13_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_10__0_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_10__1_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_10__2_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_10__3_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_10__4_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_10__5_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_10__6_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_10__7_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_10__8_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_10__9_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_10__10_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_10__11_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_10__12_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_10__13_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_11__0_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_11__1_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_11__2_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_11__3_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_11__4_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_11__5_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_11__6_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_11__7_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_11__8_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_11__9_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_11__10_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_11__11_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_11__12_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_11__13_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_12__0_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_12__1_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_12__2_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_12__3_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_12__4_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_12__5_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_12__6_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_12__7_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_12__8_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_12__9_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_12__10_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_12__11_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_12__12_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_12__13_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_13__0_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_13__1_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_13__2_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_13__3_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_13__4_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_13__5_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_13__6_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_13__7_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_13__8_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_13__9_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_13__10_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_13__11_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_13__12_,
         my_filter_adder_mult_4_multiplication_mult_21_ab_13__13_,
         my_filter_adder_mult_4_multiplication_mult_21_FS_1_n71,
         my_filter_adder_mult_4_multiplication_mult_21_FS_1_n70,
         my_filter_adder_mult_4_multiplication_mult_21_FS_1_n69,
         my_filter_adder_mult_4_multiplication_mult_21_FS_1_n68,
         my_filter_adder_mult_4_multiplication_mult_21_FS_1_n67,
         my_filter_adder_mult_4_multiplication_mult_21_FS_1_n66,
         my_filter_adder_mult_4_multiplication_mult_21_FS_1_n65,
         my_filter_adder_mult_4_multiplication_mult_21_FS_1_n64,
         my_filter_adder_mult_4_multiplication_mult_21_FS_1_n63,
         my_filter_adder_mult_4_multiplication_mult_21_FS_1_n62,
         my_filter_adder_mult_4_multiplication_mult_21_FS_1_n60,
         my_filter_adder_mult_4_multiplication_mult_21_FS_1_n59,
         my_filter_adder_mult_4_multiplication_mult_21_FS_1_n58,
         my_filter_adder_mult_4_multiplication_mult_21_FS_1_n57,
         my_filter_adder_mult_4_multiplication_mult_21_FS_1_n56,
         my_filter_adder_mult_4_multiplication_mult_21_FS_1_n55,
         my_filter_adder_mult_4_multiplication_mult_21_FS_1_n54,
         my_filter_adder_mult_4_multiplication_mult_21_FS_1_n53,
         my_filter_adder_mult_4_multiplication_mult_21_FS_1_n52,
         my_filter_adder_mult_4_multiplication_mult_21_FS_1_n51,
         my_filter_adder_mult_4_multiplication_mult_21_FS_1_n50,
         my_filter_adder_mult_4_multiplication_mult_21_FS_1_n49,
         my_filter_adder_mult_4_multiplication_mult_21_FS_1_n48,
         my_filter_adder_mult_4_multiplication_mult_21_FS_1_n47,
         my_filter_adder_mult_4_multiplication_mult_21_FS_1_n46,
         my_filter_adder_mult_4_multiplication_mult_21_FS_1_n45,
         my_filter_adder_mult_4_multiplication_mult_21_FS_1_n44,
         my_filter_adder_mult_4_multiplication_mult_21_FS_1_n43,
         my_filter_adder_mult_4_multiplication_mult_21_FS_1_n42,
         my_filter_adder_mult_4_multiplication_mult_21_FS_1_n41,
         my_filter_adder_mult_4_multiplication_mult_21_FS_1_n40,
         my_filter_adder_mult_4_multiplication_mult_21_FS_1_n39,
         my_filter_adder_mult_4_multiplication_mult_21_FS_1_n38,
         my_filter_adder_mult_4_multiplication_mult_21_FS_1_n37,
         my_filter_adder_mult_4_multiplication_mult_21_FS_1_n36,
         my_filter_adder_mult_4_multiplication_mult_21_FS_1_n35,
         my_filter_adder_mult_4_multiplication_mult_21_FS_1_n34,
         my_filter_adder_mult_4_multiplication_mult_21_FS_1_n33,
         my_filter_adder_mult_4_multiplication_mult_21_FS_1_n32,
         my_filter_adder_mult_4_multiplication_mult_21_FS_1_n31,
         my_filter_adder_mult_4_multiplication_mult_21_FS_1_n30,
         my_filter_adder_mult_4_multiplication_mult_21_FS_1_n29,
         my_filter_adder_mult_4_multiplication_mult_21_FS_1_n28,
         my_filter_adder_mult_4_multiplication_mult_21_FS_1_n27,
         my_filter_adder_mult_4_multiplication_mult_21_FS_1_n26,
         my_filter_adder_mult_4_multiplication_mult_21_FS_1_n25,
         my_filter_adder_mult_4_multiplication_mult_21_FS_1_n24,
         my_filter_adder_mult_4_multiplication_mult_21_FS_1_n23,
         my_filter_adder_mult_4_multiplication_mult_21_FS_1_n22,
         my_filter_adder_mult_4_multiplication_mult_21_FS_1_n21,
         my_filter_adder_mult_4_multiplication_mult_21_FS_1_n20,
         my_filter_adder_mult_4_multiplication_mult_21_FS_1_n19,
         my_filter_adder_mult_4_multiplication_mult_21_FS_1_n18,
         my_filter_adder_mult_4_multiplication_mult_21_FS_1_n17,
         my_filter_adder_mult_4_multiplication_mult_21_FS_1_n16,
         my_filter_adder_mult_4_multiplication_mult_21_FS_1_n15,
         my_filter_adder_mult_4_multiplication_mult_21_FS_1_n14,
         my_filter_adder_mult_4_multiplication_mult_21_FS_1_n13,
         my_filter_adder_mult_4_addition_add_19_n1,
         my_filter_adder_mult_5_multiplication_mult_21_n113,
         my_filter_adder_mult_5_multiplication_mult_21_n112,
         my_filter_adder_mult_5_multiplication_mult_21_n111,
         my_filter_adder_mult_5_multiplication_mult_21_n110,
         my_filter_adder_mult_5_multiplication_mult_21_n109,
         my_filter_adder_mult_5_multiplication_mult_21_n108,
         my_filter_adder_mult_5_multiplication_mult_21_n107,
         my_filter_adder_mult_5_multiplication_mult_21_n106,
         my_filter_adder_mult_5_multiplication_mult_21_n105,
         my_filter_adder_mult_5_multiplication_mult_21_n104,
         my_filter_adder_mult_5_multiplication_mult_21_n103,
         my_filter_adder_mult_5_multiplication_mult_21_n102,
         my_filter_adder_mult_5_multiplication_mult_21_n101,
         my_filter_adder_mult_5_multiplication_mult_21_n100,
         my_filter_adder_mult_5_multiplication_mult_21_n99,
         my_filter_adder_mult_5_multiplication_mult_21_n98,
         my_filter_adder_mult_5_multiplication_mult_21_n97,
         my_filter_adder_mult_5_multiplication_mult_21_n96,
         my_filter_adder_mult_5_multiplication_mult_21_n95,
         my_filter_adder_mult_5_multiplication_mult_21_n94,
         my_filter_adder_mult_5_multiplication_mult_21_n93,
         my_filter_adder_mult_5_multiplication_mult_21_n92,
         my_filter_adder_mult_5_multiplication_mult_21_n91,
         my_filter_adder_mult_5_multiplication_mult_21_n90,
         my_filter_adder_mult_5_multiplication_mult_21_n89,
         my_filter_adder_mult_5_multiplication_mult_21_n88,
         my_filter_adder_mult_5_multiplication_mult_21_n87,
         my_filter_adder_mult_5_multiplication_mult_21_n86,
         my_filter_adder_mult_5_multiplication_mult_21_n85,
         my_filter_adder_mult_5_multiplication_mult_21_n52,
         my_filter_adder_mult_5_multiplication_mult_21_n51,
         my_filter_adder_mult_5_multiplication_mult_21_n50,
         my_filter_adder_mult_5_multiplication_mult_21_n49,
         my_filter_adder_mult_5_multiplication_mult_21_n48,
         my_filter_adder_mult_5_multiplication_mult_21_n47,
         my_filter_adder_mult_5_multiplication_mult_21_n46,
         my_filter_adder_mult_5_multiplication_mult_21_n45,
         my_filter_adder_mult_5_multiplication_mult_21_n44,
         my_filter_adder_mult_5_multiplication_mult_21_n43,
         my_filter_adder_mult_5_multiplication_mult_21_n42,
         my_filter_adder_mult_5_multiplication_mult_21_n41,
         my_filter_adder_mult_5_multiplication_mult_21_n40,
         my_filter_adder_mult_5_multiplication_mult_21_n39,
         my_filter_adder_mult_5_multiplication_mult_21_n38,
         my_filter_adder_mult_5_multiplication_mult_21_n37,
         my_filter_adder_mult_5_multiplication_mult_21_n36,
         my_filter_adder_mult_5_multiplication_mult_21_n35,
         my_filter_adder_mult_5_multiplication_mult_21_n34,
         my_filter_adder_mult_5_multiplication_mult_21_n33,
         my_filter_adder_mult_5_multiplication_mult_21_n32,
         my_filter_adder_mult_5_multiplication_mult_21_n31,
         my_filter_adder_mult_5_multiplication_mult_21_n30,
         my_filter_adder_mult_5_multiplication_mult_21_n29,
         my_filter_adder_mult_5_multiplication_mult_21_n28,
         my_filter_adder_mult_5_multiplication_mult_21_n27,
         my_filter_adder_mult_5_multiplication_mult_21_n26,
         my_filter_adder_mult_5_multiplication_mult_21_n25,
         my_filter_adder_mult_5_multiplication_mult_21_n24,
         my_filter_adder_mult_5_multiplication_mult_21_n23,
         my_filter_adder_mult_5_multiplication_mult_21_n22,
         my_filter_adder_mult_5_multiplication_mult_21_n21,
         my_filter_adder_mult_5_multiplication_mult_21_n20,
         my_filter_adder_mult_5_multiplication_mult_21_n19,
         my_filter_adder_mult_5_multiplication_mult_21_n18,
         my_filter_adder_mult_5_multiplication_mult_21_n17,
         my_filter_adder_mult_5_multiplication_mult_21_n16,
         my_filter_adder_mult_5_multiplication_mult_21_n15,
         my_filter_adder_mult_5_multiplication_mult_21_n14,
         my_filter_adder_mult_5_multiplication_mult_21_n13,
         my_filter_adder_mult_5_multiplication_mult_21_n12,
         my_filter_adder_mult_5_multiplication_mult_21_n11,
         my_filter_adder_mult_5_multiplication_mult_21_n10,
         my_filter_adder_mult_5_multiplication_mult_21_n9,
         my_filter_adder_mult_5_multiplication_mult_21_n8,
         my_filter_adder_mult_5_multiplication_mult_21_n7,
         my_filter_adder_mult_5_multiplication_mult_21_n6,
         my_filter_adder_mult_5_multiplication_mult_21_n5,
         my_filter_adder_mult_5_multiplication_mult_21_n4,
         my_filter_adder_mult_5_multiplication_mult_21_n3,
         my_filter_adder_mult_5_multiplication_mult_21_A2_12_,
         my_filter_adder_mult_5_multiplication_mult_21_A1_0_,
         my_filter_adder_mult_5_multiplication_mult_21_A1_1_,
         my_filter_adder_mult_5_multiplication_mult_21_A1_2_,
         my_filter_adder_mult_5_multiplication_mult_21_A1_3_,
         my_filter_adder_mult_5_multiplication_mult_21_A1_4_,
         my_filter_adder_mult_5_multiplication_mult_21_A1_5_,
         my_filter_adder_mult_5_multiplication_mult_21_A1_6_,
         my_filter_adder_mult_5_multiplication_mult_21_A1_7_,
         my_filter_adder_mult_5_multiplication_mult_21_A1_8_,
         my_filter_adder_mult_5_multiplication_mult_21_A1_9_,
         my_filter_adder_mult_5_multiplication_mult_21_A1_10_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_2__1_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_2__2_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_2__3_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_2__4_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_2__5_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_2__6_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_2__7_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_2__8_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_2__9_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_2__10_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_2__11_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_2__12_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_3__1_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_3__2_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_3__3_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_3__4_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_3__5_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_3__6_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_3__7_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_3__8_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_3__9_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_3__10_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_3__11_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_3__12_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_4__1_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_4__2_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_4__3_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_4__4_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_4__5_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_4__6_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_4__7_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_4__8_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_4__9_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_4__10_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_4__11_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_4__12_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_5__1_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_5__2_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_5__3_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_5__4_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_5__5_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_5__6_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_5__7_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_5__8_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_5__9_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_5__10_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_5__11_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_5__12_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_6__1_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_6__2_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_6__3_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_6__4_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_6__5_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_6__6_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_6__7_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_6__8_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_6__9_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_6__10_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_6__11_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_6__12_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_7__1_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_7__2_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_7__3_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_7__4_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_7__5_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_7__6_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_7__7_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_7__8_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_7__9_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_7__10_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_7__11_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_7__12_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_8__1_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_8__2_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_8__3_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_8__4_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_8__5_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_8__6_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_8__7_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_8__8_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_8__9_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_8__10_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_8__11_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_8__12_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_9__1_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_9__2_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_9__3_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_9__4_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_9__5_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_9__6_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_9__7_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_9__8_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_9__9_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_9__10_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_9__11_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_9__12_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_10__1_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_10__2_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_10__3_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_10__4_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_10__5_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_10__6_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_10__7_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_10__8_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_10__9_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_10__10_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_10__11_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_10__12_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_11__1_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_11__2_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_11__3_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_11__4_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_11__5_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_11__6_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_11__7_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_11__8_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_11__9_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_11__10_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_11__11_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_11__12_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_12__1_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_12__2_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_12__3_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_12__4_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_12__5_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_12__6_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_12__7_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_12__8_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_12__9_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_12__10_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_12__11_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_12__12_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_13__0_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_13__1_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_13__2_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_13__3_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_13__4_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_13__5_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_13__6_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_13__7_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_13__8_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_13__9_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_13__10_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_13__11_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_13__12_,
         my_filter_adder_mult_5_multiplication_mult_21_SUMB_13__13_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_1__0_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_2__0_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_2__1_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_2__2_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_2__3_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_2__4_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_2__5_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_2__6_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_2__7_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_2__8_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_2__9_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_2__10_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_2__11_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_2__12_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_3__0_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_3__1_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_3__2_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_3__3_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_3__4_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_3__5_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_3__6_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_3__7_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_3__8_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_3__9_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_3__10_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_3__11_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_3__12_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_4__0_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_4__1_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_4__2_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_4__3_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_4__4_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_4__5_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_4__6_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_4__7_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_4__8_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_4__9_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_4__10_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_4__11_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_4__12_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_5__0_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_5__1_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_5__2_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_5__3_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_5__4_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_5__5_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_5__6_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_5__7_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_5__8_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_5__9_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_5__10_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_5__11_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_5__12_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_6__0_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_6__1_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_6__2_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_6__3_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_6__4_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_6__5_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_6__6_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_6__7_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_6__8_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_6__9_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_6__10_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_6__11_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_6__12_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_7__0_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_7__1_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_7__2_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_7__3_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_7__4_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_7__5_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_7__6_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_7__7_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_7__8_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_7__9_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_7__10_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_7__11_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_7__12_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_8__0_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_8__1_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_8__2_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_8__3_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_8__4_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_8__5_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_8__6_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_8__7_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_8__8_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_8__9_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_8__10_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_8__11_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_8__12_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_9__0_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_9__1_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_9__2_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_9__3_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_9__4_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_9__5_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_9__6_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_9__7_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_9__8_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_9__9_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_9__10_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_9__11_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_9__12_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_10__0_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_10__1_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_10__2_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_10__3_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_10__4_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_10__5_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_10__6_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_10__7_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_10__8_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_10__9_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_10__10_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_10__11_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_10__12_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_11__0_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_11__1_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_11__2_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_11__3_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_11__4_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_11__5_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_11__6_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_11__7_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_11__8_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_11__9_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_11__10_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_11__11_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_11__12_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_12__0_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_12__1_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_12__2_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_12__3_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_12__4_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_12__5_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_12__6_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_12__7_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_12__8_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_12__9_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_12__10_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_12__11_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_12__12_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_13__0_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_13__1_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_13__2_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_13__3_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_13__4_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_13__5_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_13__6_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_13__7_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_13__8_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_13__9_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_13__10_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_13__11_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_13__12_,
         my_filter_adder_mult_5_multiplication_mult_21_CARRYB_13__13_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_0__2_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_0__3_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_0__4_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_0__5_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_0__6_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_0__7_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_0__8_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_0__9_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_0__10_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_0__11_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_0__12_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_0__13_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_1__1_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_1__2_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_1__3_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_1__4_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_1__5_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_1__6_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_1__7_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_1__8_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_1__9_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_1__10_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_1__11_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_1__12_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_1__13_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_2__0_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_2__1_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_2__2_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_2__3_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_2__4_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_2__5_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_2__6_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_2__7_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_2__8_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_2__9_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_2__10_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_2__11_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_2__12_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_2__13_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_3__0_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_3__1_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_3__2_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_3__3_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_3__4_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_3__5_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_3__6_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_3__7_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_3__8_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_3__9_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_3__10_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_3__11_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_3__12_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_3__13_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_4__0_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_4__1_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_4__2_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_4__3_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_4__4_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_4__5_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_4__6_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_4__7_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_4__8_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_4__9_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_4__10_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_4__11_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_4__12_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_4__13_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_5__0_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_5__1_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_5__2_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_5__3_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_5__4_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_5__5_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_5__6_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_5__7_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_5__8_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_5__9_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_5__10_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_5__11_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_5__12_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_5__13_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_6__0_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_6__1_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_6__2_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_6__3_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_6__4_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_6__5_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_6__6_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_6__7_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_6__8_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_6__9_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_6__10_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_6__11_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_6__12_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_6__13_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_7__0_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_7__1_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_7__2_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_7__3_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_7__4_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_7__5_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_7__6_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_7__7_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_7__8_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_7__9_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_7__10_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_7__11_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_7__12_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_7__13_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_8__0_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_8__1_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_8__2_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_8__3_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_8__4_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_8__5_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_8__6_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_8__7_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_8__8_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_8__9_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_8__10_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_8__11_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_8__12_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_8__13_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_9__0_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_9__1_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_9__2_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_9__3_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_9__4_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_9__5_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_9__6_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_9__7_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_9__8_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_9__9_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_9__10_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_9__11_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_9__12_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_9__13_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_10__0_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_10__1_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_10__2_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_10__3_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_10__4_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_10__5_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_10__6_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_10__7_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_10__8_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_10__9_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_10__10_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_10__11_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_10__12_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_10__13_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_11__0_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_11__1_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_11__2_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_11__3_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_11__4_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_11__5_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_11__6_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_11__7_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_11__8_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_11__9_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_11__10_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_11__11_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_11__12_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_11__13_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_12__0_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_12__1_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_12__2_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_12__3_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_12__4_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_12__5_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_12__6_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_12__7_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_12__8_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_12__9_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_12__10_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_12__11_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_12__12_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_12__13_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_13__0_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_13__1_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_13__2_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_13__3_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_13__4_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_13__5_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_13__6_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_13__7_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_13__8_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_13__9_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_13__10_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_13__11_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_13__12_,
         my_filter_adder_mult_5_multiplication_mult_21_ab_13__13_,
         my_filter_adder_mult_5_multiplication_mult_21_FS_1_n71,
         my_filter_adder_mult_5_multiplication_mult_21_FS_1_n70,
         my_filter_adder_mult_5_multiplication_mult_21_FS_1_n69,
         my_filter_adder_mult_5_multiplication_mult_21_FS_1_n68,
         my_filter_adder_mult_5_multiplication_mult_21_FS_1_n67,
         my_filter_adder_mult_5_multiplication_mult_21_FS_1_n66,
         my_filter_adder_mult_5_multiplication_mult_21_FS_1_n65,
         my_filter_adder_mult_5_multiplication_mult_21_FS_1_n64,
         my_filter_adder_mult_5_multiplication_mult_21_FS_1_n63,
         my_filter_adder_mult_5_multiplication_mult_21_FS_1_n62,
         my_filter_adder_mult_5_multiplication_mult_21_FS_1_n60,
         my_filter_adder_mult_5_multiplication_mult_21_FS_1_n59,
         my_filter_adder_mult_5_multiplication_mult_21_FS_1_n58,
         my_filter_adder_mult_5_multiplication_mult_21_FS_1_n57,
         my_filter_adder_mult_5_multiplication_mult_21_FS_1_n56,
         my_filter_adder_mult_5_multiplication_mult_21_FS_1_n55,
         my_filter_adder_mult_5_multiplication_mult_21_FS_1_n54,
         my_filter_adder_mult_5_multiplication_mult_21_FS_1_n53,
         my_filter_adder_mult_5_multiplication_mult_21_FS_1_n52,
         my_filter_adder_mult_5_multiplication_mult_21_FS_1_n51,
         my_filter_adder_mult_5_multiplication_mult_21_FS_1_n50,
         my_filter_adder_mult_5_multiplication_mult_21_FS_1_n49,
         my_filter_adder_mult_5_multiplication_mult_21_FS_1_n48,
         my_filter_adder_mult_5_multiplication_mult_21_FS_1_n47,
         my_filter_adder_mult_5_multiplication_mult_21_FS_1_n46,
         my_filter_adder_mult_5_multiplication_mult_21_FS_1_n45,
         my_filter_adder_mult_5_multiplication_mult_21_FS_1_n44,
         my_filter_adder_mult_5_multiplication_mult_21_FS_1_n43,
         my_filter_adder_mult_5_multiplication_mult_21_FS_1_n42,
         my_filter_adder_mult_5_multiplication_mult_21_FS_1_n41,
         my_filter_adder_mult_5_multiplication_mult_21_FS_1_n40,
         my_filter_adder_mult_5_multiplication_mult_21_FS_1_n39,
         my_filter_adder_mult_5_multiplication_mult_21_FS_1_n38,
         my_filter_adder_mult_5_multiplication_mult_21_FS_1_n37,
         my_filter_adder_mult_5_multiplication_mult_21_FS_1_n36,
         my_filter_adder_mult_5_multiplication_mult_21_FS_1_n35,
         my_filter_adder_mult_5_multiplication_mult_21_FS_1_n34,
         my_filter_adder_mult_5_multiplication_mult_21_FS_1_n33,
         my_filter_adder_mult_5_multiplication_mult_21_FS_1_n32,
         my_filter_adder_mult_5_multiplication_mult_21_FS_1_n31,
         my_filter_adder_mult_5_multiplication_mult_21_FS_1_n30,
         my_filter_adder_mult_5_multiplication_mult_21_FS_1_n29,
         my_filter_adder_mult_5_multiplication_mult_21_FS_1_n28,
         my_filter_adder_mult_5_multiplication_mult_21_FS_1_n27,
         my_filter_adder_mult_5_multiplication_mult_21_FS_1_n26,
         my_filter_adder_mult_5_multiplication_mult_21_FS_1_n25,
         my_filter_adder_mult_5_multiplication_mult_21_FS_1_n24,
         my_filter_adder_mult_5_multiplication_mult_21_FS_1_n23,
         my_filter_adder_mult_5_multiplication_mult_21_FS_1_n22,
         my_filter_adder_mult_5_multiplication_mult_21_FS_1_n21,
         my_filter_adder_mult_5_multiplication_mult_21_FS_1_n20,
         my_filter_adder_mult_5_multiplication_mult_21_FS_1_n19,
         my_filter_adder_mult_5_multiplication_mult_21_FS_1_n18,
         my_filter_adder_mult_5_multiplication_mult_21_FS_1_n17,
         my_filter_adder_mult_5_multiplication_mult_21_FS_1_n16,
         my_filter_adder_mult_5_multiplication_mult_21_FS_1_n15,
         my_filter_adder_mult_5_multiplication_mult_21_FS_1_n14,
         my_filter_adder_mult_5_multiplication_mult_21_FS_1_n13,
         my_filter_adder_mult_5_addition_add_19_n1,
         my_filter_adder_mult_6_multiplication_mult_21_n113,
         my_filter_adder_mult_6_multiplication_mult_21_n112,
         my_filter_adder_mult_6_multiplication_mult_21_n111,
         my_filter_adder_mult_6_multiplication_mult_21_n110,
         my_filter_adder_mult_6_multiplication_mult_21_n109,
         my_filter_adder_mult_6_multiplication_mult_21_n108,
         my_filter_adder_mult_6_multiplication_mult_21_n107,
         my_filter_adder_mult_6_multiplication_mult_21_n106,
         my_filter_adder_mult_6_multiplication_mult_21_n105,
         my_filter_adder_mult_6_multiplication_mult_21_n104,
         my_filter_adder_mult_6_multiplication_mult_21_n103,
         my_filter_adder_mult_6_multiplication_mult_21_n102,
         my_filter_adder_mult_6_multiplication_mult_21_n101,
         my_filter_adder_mult_6_multiplication_mult_21_n100,
         my_filter_adder_mult_6_multiplication_mult_21_n99,
         my_filter_adder_mult_6_multiplication_mult_21_n98,
         my_filter_adder_mult_6_multiplication_mult_21_n97,
         my_filter_adder_mult_6_multiplication_mult_21_n96,
         my_filter_adder_mult_6_multiplication_mult_21_n95,
         my_filter_adder_mult_6_multiplication_mult_21_n94,
         my_filter_adder_mult_6_multiplication_mult_21_n93,
         my_filter_adder_mult_6_multiplication_mult_21_n92,
         my_filter_adder_mult_6_multiplication_mult_21_n91,
         my_filter_adder_mult_6_multiplication_mult_21_n90,
         my_filter_adder_mult_6_multiplication_mult_21_n89,
         my_filter_adder_mult_6_multiplication_mult_21_n88,
         my_filter_adder_mult_6_multiplication_mult_21_n87,
         my_filter_adder_mult_6_multiplication_mult_21_n86,
         my_filter_adder_mult_6_multiplication_mult_21_n85,
         my_filter_adder_mult_6_multiplication_mult_21_n52,
         my_filter_adder_mult_6_multiplication_mult_21_n51,
         my_filter_adder_mult_6_multiplication_mult_21_n50,
         my_filter_adder_mult_6_multiplication_mult_21_n49,
         my_filter_adder_mult_6_multiplication_mult_21_n48,
         my_filter_adder_mult_6_multiplication_mult_21_n47,
         my_filter_adder_mult_6_multiplication_mult_21_n46,
         my_filter_adder_mult_6_multiplication_mult_21_n45,
         my_filter_adder_mult_6_multiplication_mult_21_n44,
         my_filter_adder_mult_6_multiplication_mult_21_n43,
         my_filter_adder_mult_6_multiplication_mult_21_n42,
         my_filter_adder_mult_6_multiplication_mult_21_n41,
         my_filter_adder_mult_6_multiplication_mult_21_n40,
         my_filter_adder_mult_6_multiplication_mult_21_n39,
         my_filter_adder_mult_6_multiplication_mult_21_n38,
         my_filter_adder_mult_6_multiplication_mult_21_n37,
         my_filter_adder_mult_6_multiplication_mult_21_n36,
         my_filter_adder_mult_6_multiplication_mult_21_n35,
         my_filter_adder_mult_6_multiplication_mult_21_n34,
         my_filter_adder_mult_6_multiplication_mult_21_n33,
         my_filter_adder_mult_6_multiplication_mult_21_n32,
         my_filter_adder_mult_6_multiplication_mult_21_n31,
         my_filter_adder_mult_6_multiplication_mult_21_n30,
         my_filter_adder_mult_6_multiplication_mult_21_n29,
         my_filter_adder_mult_6_multiplication_mult_21_n28,
         my_filter_adder_mult_6_multiplication_mult_21_n27,
         my_filter_adder_mult_6_multiplication_mult_21_n26,
         my_filter_adder_mult_6_multiplication_mult_21_n25,
         my_filter_adder_mult_6_multiplication_mult_21_n24,
         my_filter_adder_mult_6_multiplication_mult_21_n23,
         my_filter_adder_mult_6_multiplication_mult_21_n22,
         my_filter_adder_mult_6_multiplication_mult_21_n21,
         my_filter_adder_mult_6_multiplication_mult_21_n20,
         my_filter_adder_mult_6_multiplication_mult_21_n19,
         my_filter_adder_mult_6_multiplication_mult_21_n18,
         my_filter_adder_mult_6_multiplication_mult_21_n17,
         my_filter_adder_mult_6_multiplication_mult_21_n16,
         my_filter_adder_mult_6_multiplication_mult_21_n15,
         my_filter_adder_mult_6_multiplication_mult_21_n14,
         my_filter_adder_mult_6_multiplication_mult_21_n13,
         my_filter_adder_mult_6_multiplication_mult_21_n12,
         my_filter_adder_mult_6_multiplication_mult_21_n11,
         my_filter_adder_mult_6_multiplication_mult_21_n10,
         my_filter_adder_mult_6_multiplication_mult_21_n9,
         my_filter_adder_mult_6_multiplication_mult_21_n8,
         my_filter_adder_mult_6_multiplication_mult_21_n7,
         my_filter_adder_mult_6_multiplication_mult_21_n6,
         my_filter_adder_mult_6_multiplication_mult_21_n5,
         my_filter_adder_mult_6_multiplication_mult_21_n4,
         my_filter_adder_mult_6_multiplication_mult_21_n3,
         my_filter_adder_mult_6_multiplication_mult_21_A2_12_,
         my_filter_adder_mult_6_multiplication_mult_21_A1_0_,
         my_filter_adder_mult_6_multiplication_mult_21_A1_1_,
         my_filter_adder_mult_6_multiplication_mult_21_A1_2_,
         my_filter_adder_mult_6_multiplication_mult_21_A1_3_,
         my_filter_adder_mult_6_multiplication_mult_21_A1_4_,
         my_filter_adder_mult_6_multiplication_mult_21_A1_5_,
         my_filter_adder_mult_6_multiplication_mult_21_A1_6_,
         my_filter_adder_mult_6_multiplication_mult_21_A1_7_,
         my_filter_adder_mult_6_multiplication_mult_21_A1_8_,
         my_filter_adder_mult_6_multiplication_mult_21_A1_9_,
         my_filter_adder_mult_6_multiplication_mult_21_A1_10_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_2__1_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_2__2_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_2__3_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_2__4_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_2__5_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_2__6_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_2__7_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_2__8_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_2__9_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_2__10_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_2__11_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_2__12_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_3__1_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_3__2_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_3__3_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_3__4_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_3__5_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_3__6_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_3__7_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_3__8_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_3__9_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_3__10_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_3__11_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_3__12_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_4__1_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_4__2_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_4__3_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_4__4_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_4__5_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_4__6_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_4__7_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_4__8_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_4__9_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_4__10_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_4__11_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_4__12_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_5__1_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_5__2_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_5__3_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_5__4_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_5__5_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_5__6_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_5__7_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_5__8_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_5__9_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_5__10_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_5__11_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_5__12_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_6__1_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_6__2_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_6__3_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_6__4_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_6__5_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_6__6_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_6__7_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_6__8_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_6__9_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_6__10_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_6__11_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_6__12_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_7__1_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_7__2_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_7__3_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_7__4_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_7__5_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_7__6_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_7__7_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_7__8_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_7__9_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_7__10_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_7__11_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_7__12_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_8__1_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_8__2_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_8__3_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_8__4_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_8__5_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_8__6_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_8__7_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_8__8_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_8__9_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_8__10_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_8__11_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_8__12_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_9__1_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_9__2_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_9__3_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_9__4_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_9__5_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_9__6_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_9__7_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_9__8_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_9__9_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_9__10_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_9__11_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_9__12_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_10__1_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_10__2_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_10__3_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_10__4_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_10__5_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_10__6_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_10__7_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_10__8_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_10__9_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_10__10_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_10__11_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_10__12_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_11__1_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_11__2_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_11__3_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_11__4_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_11__5_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_11__6_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_11__7_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_11__8_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_11__9_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_11__10_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_11__11_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_11__12_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_12__1_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_12__2_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_12__3_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_12__4_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_12__5_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_12__6_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_12__7_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_12__8_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_12__9_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_12__10_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_12__11_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_12__12_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_13__0_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_13__1_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_13__2_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_13__3_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_13__4_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_13__5_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_13__6_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_13__7_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_13__8_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_13__9_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_13__10_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_13__11_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_13__12_,
         my_filter_adder_mult_6_multiplication_mult_21_SUMB_13__13_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_1__0_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_2__0_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_2__1_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_2__2_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_2__3_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_2__4_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_2__5_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_2__6_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_2__7_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_2__8_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_2__9_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_2__10_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_2__11_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_2__12_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_3__0_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_3__1_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_3__2_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_3__3_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_3__4_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_3__5_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_3__6_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_3__7_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_3__8_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_3__9_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_3__10_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_3__11_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_3__12_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_4__0_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_4__1_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_4__2_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_4__3_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_4__4_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_4__5_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_4__6_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_4__7_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_4__8_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_4__9_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_4__10_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_4__11_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_4__12_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_5__0_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_5__1_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_5__2_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_5__3_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_5__4_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_5__5_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_5__6_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_5__7_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_5__8_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_5__9_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_5__10_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_5__11_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_5__12_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_6__0_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_6__1_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_6__2_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_6__3_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_6__4_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_6__5_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_6__6_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_6__7_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_6__8_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_6__9_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_6__10_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_6__11_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_6__12_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_7__0_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_7__1_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_7__2_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_7__3_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_7__4_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_7__5_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_7__6_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_7__7_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_7__8_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_7__9_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_7__10_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_7__11_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_7__12_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_8__0_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_8__1_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_8__2_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_8__3_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_8__4_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_8__5_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_8__6_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_8__7_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_8__8_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_8__9_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_8__10_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_8__11_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_8__12_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_9__0_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_9__1_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_9__2_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_9__3_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_9__4_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_9__5_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_9__6_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_9__7_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_9__8_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_9__9_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_9__10_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_9__11_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_9__12_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_10__0_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_10__1_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_10__2_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_10__3_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_10__4_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_10__5_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_10__6_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_10__7_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_10__8_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_10__9_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_10__10_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_10__11_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_10__12_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_11__0_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_11__1_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_11__2_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_11__3_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_11__4_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_11__5_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_11__6_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_11__7_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_11__8_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_11__9_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_11__10_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_11__11_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_11__12_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_12__0_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_12__1_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_12__2_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_12__3_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_12__4_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_12__5_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_12__6_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_12__7_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_12__8_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_12__9_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_12__10_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_12__11_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_12__12_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_13__0_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_13__1_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_13__2_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_13__3_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_13__4_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_13__5_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_13__6_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_13__7_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_13__8_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_13__9_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_13__10_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_13__11_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_13__12_,
         my_filter_adder_mult_6_multiplication_mult_21_CARRYB_13__13_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_0__2_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_0__3_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_0__4_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_0__5_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_0__6_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_0__7_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_0__8_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_0__9_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_0__10_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_0__11_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_0__12_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_0__13_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_1__1_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_1__2_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_1__3_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_1__4_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_1__5_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_1__6_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_1__7_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_1__8_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_1__9_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_1__10_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_1__11_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_1__12_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_1__13_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_2__0_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_2__1_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_2__2_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_2__3_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_2__4_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_2__5_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_2__6_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_2__7_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_2__8_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_2__9_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_2__10_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_2__11_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_2__12_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_2__13_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_3__0_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_3__1_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_3__2_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_3__3_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_3__4_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_3__5_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_3__6_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_3__7_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_3__8_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_3__9_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_3__10_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_3__11_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_3__12_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_3__13_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_4__0_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_4__1_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_4__2_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_4__3_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_4__4_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_4__5_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_4__6_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_4__7_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_4__8_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_4__9_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_4__10_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_4__11_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_4__12_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_4__13_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_5__0_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_5__1_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_5__2_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_5__3_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_5__4_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_5__5_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_5__6_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_5__7_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_5__8_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_5__9_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_5__10_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_5__11_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_5__12_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_5__13_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_6__0_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_6__1_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_6__2_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_6__3_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_6__4_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_6__5_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_6__6_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_6__7_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_6__8_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_6__9_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_6__10_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_6__11_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_6__12_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_6__13_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_7__0_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_7__1_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_7__2_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_7__3_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_7__4_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_7__5_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_7__6_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_7__7_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_7__8_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_7__9_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_7__10_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_7__11_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_7__12_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_7__13_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_8__0_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_8__1_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_8__2_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_8__3_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_8__4_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_8__5_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_8__6_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_8__7_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_8__8_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_8__9_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_8__10_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_8__11_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_8__12_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_8__13_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_9__0_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_9__1_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_9__2_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_9__3_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_9__4_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_9__5_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_9__6_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_9__7_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_9__8_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_9__9_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_9__10_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_9__11_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_9__12_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_9__13_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_10__0_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_10__1_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_10__2_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_10__3_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_10__4_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_10__5_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_10__6_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_10__7_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_10__8_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_10__9_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_10__10_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_10__11_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_10__12_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_10__13_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_11__0_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_11__1_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_11__2_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_11__3_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_11__4_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_11__5_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_11__6_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_11__7_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_11__8_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_11__9_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_11__10_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_11__11_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_11__12_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_11__13_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_12__0_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_12__1_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_12__2_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_12__3_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_12__4_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_12__5_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_12__6_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_12__7_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_12__8_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_12__9_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_12__10_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_12__11_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_12__12_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_12__13_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_13__0_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_13__1_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_13__2_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_13__3_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_13__4_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_13__5_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_13__6_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_13__7_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_13__8_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_13__9_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_13__10_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_13__11_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_13__12_,
         my_filter_adder_mult_6_multiplication_mult_21_ab_13__13_,
         my_filter_adder_mult_6_multiplication_mult_21_FS_1_n71,
         my_filter_adder_mult_6_multiplication_mult_21_FS_1_n70,
         my_filter_adder_mult_6_multiplication_mult_21_FS_1_n69,
         my_filter_adder_mult_6_multiplication_mult_21_FS_1_n68,
         my_filter_adder_mult_6_multiplication_mult_21_FS_1_n67,
         my_filter_adder_mult_6_multiplication_mult_21_FS_1_n66,
         my_filter_adder_mult_6_multiplication_mult_21_FS_1_n65,
         my_filter_adder_mult_6_multiplication_mult_21_FS_1_n64,
         my_filter_adder_mult_6_multiplication_mult_21_FS_1_n63,
         my_filter_adder_mult_6_multiplication_mult_21_FS_1_n62,
         my_filter_adder_mult_6_multiplication_mult_21_FS_1_n60,
         my_filter_adder_mult_6_multiplication_mult_21_FS_1_n59,
         my_filter_adder_mult_6_multiplication_mult_21_FS_1_n58,
         my_filter_adder_mult_6_multiplication_mult_21_FS_1_n57,
         my_filter_adder_mult_6_multiplication_mult_21_FS_1_n56,
         my_filter_adder_mult_6_multiplication_mult_21_FS_1_n55,
         my_filter_adder_mult_6_multiplication_mult_21_FS_1_n54,
         my_filter_adder_mult_6_multiplication_mult_21_FS_1_n53,
         my_filter_adder_mult_6_multiplication_mult_21_FS_1_n52,
         my_filter_adder_mult_6_multiplication_mult_21_FS_1_n51,
         my_filter_adder_mult_6_multiplication_mult_21_FS_1_n50,
         my_filter_adder_mult_6_multiplication_mult_21_FS_1_n49,
         my_filter_adder_mult_6_multiplication_mult_21_FS_1_n48,
         my_filter_adder_mult_6_multiplication_mult_21_FS_1_n47,
         my_filter_adder_mult_6_multiplication_mult_21_FS_1_n46,
         my_filter_adder_mult_6_multiplication_mult_21_FS_1_n45,
         my_filter_adder_mult_6_multiplication_mult_21_FS_1_n44,
         my_filter_adder_mult_6_multiplication_mult_21_FS_1_n43,
         my_filter_adder_mult_6_multiplication_mult_21_FS_1_n42,
         my_filter_adder_mult_6_multiplication_mult_21_FS_1_n41,
         my_filter_adder_mult_6_multiplication_mult_21_FS_1_n40,
         my_filter_adder_mult_6_multiplication_mult_21_FS_1_n39,
         my_filter_adder_mult_6_multiplication_mult_21_FS_1_n38,
         my_filter_adder_mult_6_multiplication_mult_21_FS_1_n37,
         my_filter_adder_mult_6_multiplication_mult_21_FS_1_n36,
         my_filter_adder_mult_6_multiplication_mult_21_FS_1_n35,
         my_filter_adder_mult_6_multiplication_mult_21_FS_1_n34,
         my_filter_adder_mult_6_multiplication_mult_21_FS_1_n33,
         my_filter_adder_mult_6_multiplication_mult_21_FS_1_n32,
         my_filter_adder_mult_6_multiplication_mult_21_FS_1_n31,
         my_filter_adder_mult_6_multiplication_mult_21_FS_1_n30,
         my_filter_adder_mult_6_multiplication_mult_21_FS_1_n29,
         my_filter_adder_mult_6_multiplication_mult_21_FS_1_n28,
         my_filter_adder_mult_6_multiplication_mult_21_FS_1_n27,
         my_filter_adder_mult_6_multiplication_mult_21_FS_1_n26,
         my_filter_adder_mult_6_multiplication_mult_21_FS_1_n25,
         my_filter_adder_mult_6_multiplication_mult_21_FS_1_n24,
         my_filter_adder_mult_6_multiplication_mult_21_FS_1_n23,
         my_filter_adder_mult_6_multiplication_mult_21_FS_1_n22,
         my_filter_adder_mult_6_multiplication_mult_21_FS_1_n21,
         my_filter_adder_mult_6_multiplication_mult_21_FS_1_n20,
         my_filter_adder_mult_6_multiplication_mult_21_FS_1_n19,
         my_filter_adder_mult_6_multiplication_mult_21_FS_1_n18,
         my_filter_adder_mult_6_multiplication_mult_21_FS_1_n17,
         my_filter_adder_mult_6_multiplication_mult_21_FS_1_n16,
         my_filter_adder_mult_6_multiplication_mult_21_FS_1_n15,
         my_filter_adder_mult_6_multiplication_mult_21_FS_1_n14,
         my_filter_adder_mult_6_multiplication_mult_21_FS_1_n13,
         my_filter_adder_mult_6_addition_add_19_n1,
         my_filter_adder_mult_7_multiplication_mult_21_n113,
         my_filter_adder_mult_7_multiplication_mult_21_n112,
         my_filter_adder_mult_7_multiplication_mult_21_n111,
         my_filter_adder_mult_7_multiplication_mult_21_n110,
         my_filter_adder_mult_7_multiplication_mult_21_n109,
         my_filter_adder_mult_7_multiplication_mult_21_n108,
         my_filter_adder_mult_7_multiplication_mult_21_n107,
         my_filter_adder_mult_7_multiplication_mult_21_n106,
         my_filter_adder_mult_7_multiplication_mult_21_n105,
         my_filter_adder_mult_7_multiplication_mult_21_n104,
         my_filter_adder_mult_7_multiplication_mult_21_n103,
         my_filter_adder_mult_7_multiplication_mult_21_n102,
         my_filter_adder_mult_7_multiplication_mult_21_n101,
         my_filter_adder_mult_7_multiplication_mult_21_n100,
         my_filter_adder_mult_7_multiplication_mult_21_n99,
         my_filter_adder_mult_7_multiplication_mult_21_n98,
         my_filter_adder_mult_7_multiplication_mult_21_n97,
         my_filter_adder_mult_7_multiplication_mult_21_n96,
         my_filter_adder_mult_7_multiplication_mult_21_n95,
         my_filter_adder_mult_7_multiplication_mult_21_n94,
         my_filter_adder_mult_7_multiplication_mult_21_n93,
         my_filter_adder_mult_7_multiplication_mult_21_n92,
         my_filter_adder_mult_7_multiplication_mult_21_n91,
         my_filter_adder_mult_7_multiplication_mult_21_n90,
         my_filter_adder_mult_7_multiplication_mult_21_n89,
         my_filter_adder_mult_7_multiplication_mult_21_n88,
         my_filter_adder_mult_7_multiplication_mult_21_n87,
         my_filter_adder_mult_7_multiplication_mult_21_n86,
         my_filter_adder_mult_7_multiplication_mult_21_n85,
         my_filter_adder_mult_7_multiplication_mult_21_n52,
         my_filter_adder_mult_7_multiplication_mult_21_n51,
         my_filter_adder_mult_7_multiplication_mult_21_n50,
         my_filter_adder_mult_7_multiplication_mult_21_n49,
         my_filter_adder_mult_7_multiplication_mult_21_n48,
         my_filter_adder_mult_7_multiplication_mult_21_n47,
         my_filter_adder_mult_7_multiplication_mult_21_n46,
         my_filter_adder_mult_7_multiplication_mult_21_n45,
         my_filter_adder_mult_7_multiplication_mult_21_n44,
         my_filter_adder_mult_7_multiplication_mult_21_n43,
         my_filter_adder_mult_7_multiplication_mult_21_n42,
         my_filter_adder_mult_7_multiplication_mult_21_n41,
         my_filter_adder_mult_7_multiplication_mult_21_n40,
         my_filter_adder_mult_7_multiplication_mult_21_n39,
         my_filter_adder_mult_7_multiplication_mult_21_n38,
         my_filter_adder_mult_7_multiplication_mult_21_n37,
         my_filter_adder_mult_7_multiplication_mult_21_n36,
         my_filter_adder_mult_7_multiplication_mult_21_n35,
         my_filter_adder_mult_7_multiplication_mult_21_n34,
         my_filter_adder_mult_7_multiplication_mult_21_n33,
         my_filter_adder_mult_7_multiplication_mult_21_n32,
         my_filter_adder_mult_7_multiplication_mult_21_n31,
         my_filter_adder_mult_7_multiplication_mult_21_n30,
         my_filter_adder_mult_7_multiplication_mult_21_n29,
         my_filter_adder_mult_7_multiplication_mult_21_n28,
         my_filter_adder_mult_7_multiplication_mult_21_n27,
         my_filter_adder_mult_7_multiplication_mult_21_n26,
         my_filter_adder_mult_7_multiplication_mult_21_n25,
         my_filter_adder_mult_7_multiplication_mult_21_n24,
         my_filter_adder_mult_7_multiplication_mult_21_n23,
         my_filter_adder_mult_7_multiplication_mult_21_n22,
         my_filter_adder_mult_7_multiplication_mult_21_n21,
         my_filter_adder_mult_7_multiplication_mult_21_n20,
         my_filter_adder_mult_7_multiplication_mult_21_n19,
         my_filter_adder_mult_7_multiplication_mult_21_n18,
         my_filter_adder_mult_7_multiplication_mult_21_n17,
         my_filter_adder_mult_7_multiplication_mult_21_n16,
         my_filter_adder_mult_7_multiplication_mult_21_n15,
         my_filter_adder_mult_7_multiplication_mult_21_n14,
         my_filter_adder_mult_7_multiplication_mult_21_n13,
         my_filter_adder_mult_7_multiplication_mult_21_n12,
         my_filter_adder_mult_7_multiplication_mult_21_n11,
         my_filter_adder_mult_7_multiplication_mult_21_n10,
         my_filter_adder_mult_7_multiplication_mult_21_n9,
         my_filter_adder_mult_7_multiplication_mult_21_n8,
         my_filter_adder_mult_7_multiplication_mult_21_n7,
         my_filter_adder_mult_7_multiplication_mult_21_n6,
         my_filter_adder_mult_7_multiplication_mult_21_n5,
         my_filter_adder_mult_7_multiplication_mult_21_n4,
         my_filter_adder_mult_7_multiplication_mult_21_n3,
         my_filter_adder_mult_7_multiplication_mult_21_A2_12_,
         my_filter_adder_mult_7_multiplication_mult_21_A1_0_,
         my_filter_adder_mult_7_multiplication_mult_21_A1_1_,
         my_filter_adder_mult_7_multiplication_mult_21_A1_2_,
         my_filter_adder_mult_7_multiplication_mult_21_A1_3_,
         my_filter_adder_mult_7_multiplication_mult_21_A1_4_,
         my_filter_adder_mult_7_multiplication_mult_21_A1_5_,
         my_filter_adder_mult_7_multiplication_mult_21_A1_6_,
         my_filter_adder_mult_7_multiplication_mult_21_A1_7_,
         my_filter_adder_mult_7_multiplication_mult_21_A1_8_,
         my_filter_adder_mult_7_multiplication_mult_21_A1_9_,
         my_filter_adder_mult_7_multiplication_mult_21_A1_10_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_2__1_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_2__2_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_2__3_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_2__4_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_2__5_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_2__6_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_2__7_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_2__8_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_2__9_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_2__10_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_2__11_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_2__12_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_3__1_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_3__2_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_3__3_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_3__4_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_3__5_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_3__6_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_3__7_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_3__8_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_3__9_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_3__10_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_3__11_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_3__12_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_4__1_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_4__2_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_4__3_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_4__4_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_4__5_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_4__6_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_4__7_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_4__8_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_4__9_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_4__10_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_4__11_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_4__12_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_5__1_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_5__2_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_5__3_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_5__4_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_5__5_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_5__6_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_5__7_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_5__8_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_5__9_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_5__10_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_5__11_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_5__12_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_6__1_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_6__2_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_6__3_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_6__4_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_6__5_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_6__6_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_6__7_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_6__8_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_6__9_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_6__10_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_6__11_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_6__12_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_7__1_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_7__2_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_7__3_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_7__4_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_7__5_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_7__6_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_7__7_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_7__8_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_7__9_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_7__10_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_7__11_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_7__12_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_8__1_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_8__2_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_8__3_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_8__4_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_8__5_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_8__6_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_8__7_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_8__8_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_8__9_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_8__10_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_8__11_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_8__12_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_9__1_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_9__2_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_9__3_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_9__4_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_9__5_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_9__6_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_9__7_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_9__8_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_9__9_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_9__10_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_9__11_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_9__12_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_10__1_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_10__2_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_10__3_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_10__4_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_10__5_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_10__6_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_10__7_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_10__8_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_10__9_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_10__10_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_10__11_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_10__12_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_11__1_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_11__2_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_11__3_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_11__4_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_11__5_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_11__6_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_11__7_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_11__8_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_11__9_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_11__10_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_11__11_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_11__12_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_12__1_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_12__2_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_12__3_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_12__4_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_12__5_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_12__6_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_12__7_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_12__8_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_12__9_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_12__10_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_12__11_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_12__12_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_13__0_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_13__1_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_13__2_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_13__3_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_13__4_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_13__5_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_13__6_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_13__7_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_13__8_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_13__9_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_13__10_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_13__11_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_13__12_,
         my_filter_adder_mult_7_multiplication_mult_21_SUMB_13__13_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_1__0_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_2__0_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_2__1_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_2__2_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_2__3_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_2__4_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_2__5_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_2__6_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_2__7_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_2__8_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_2__9_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_2__10_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_2__11_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_2__12_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_3__0_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_3__1_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_3__2_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_3__3_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_3__4_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_3__5_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_3__6_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_3__7_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_3__8_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_3__9_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_3__10_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_3__11_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_3__12_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_4__0_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_4__1_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_4__2_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_4__3_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_4__4_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_4__5_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_4__6_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_4__7_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_4__8_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_4__9_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_4__10_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_4__11_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_4__12_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_5__0_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_5__1_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_5__2_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_5__3_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_5__4_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_5__5_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_5__6_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_5__7_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_5__8_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_5__9_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_5__10_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_5__11_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_5__12_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_6__0_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_6__1_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_6__2_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_6__3_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_6__4_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_6__5_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_6__6_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_6__7_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_6__8_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_6__9_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_6__10_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_6__11_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_6__12_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_7__0_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_7__1_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_7__2_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_7__3_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_7__4_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_7__5_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_7__6_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_7__7_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_7__8_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_7__9_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_7__10_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_7__11_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_7__12_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_8__0_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_8__1_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_8__2_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_8__3_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_8__4_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_8__5_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_8__6_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_8__7_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_8__8_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_8__9_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_8__10_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_8__11_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_8__12_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_9__0_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_9__1_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_9__2_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_9__3_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_9__4_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_9__5_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_9__6_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_9__7_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_9__8_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_9__9_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_9__10_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_9__11_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_9__12_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_10__0_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_10__1_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_10__2_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_10__3_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_10__4_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_10__5_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_10__6_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_10__7_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_10__8_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_10__9_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_10__10_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_10__11_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_10__12_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_11__0_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_11__1_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_11__2_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_11__3_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_11__4_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_11__5_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_11__6_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_11__7_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_11__8_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_11__9_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_11__10_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_11__11_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_11__12_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_12__0_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_12__1_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_12__2_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_12__3_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_12__4_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_12__5_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_12__6_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_12__7_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_12__8_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_12__9_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_12__10_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_12__11_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_12__12_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_13__0_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_13__1_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_13__2_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_13__3_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_13__4_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_13__5_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_13__6_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_13__7_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_13__8_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_13__9_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_13__10_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_13__11_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_13__12_,
         my_filter_adder_mult_7_multiplication_mult_21_CARRYB_13__13_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_0__2_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_0__3_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_0__4_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_0__5_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_0__6_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_0__7_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_0__8_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_0__9_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_0__10_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_0__11_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_0__12_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_0__13_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_1__1_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_1__2_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_1__3_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_1__4_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_1__5_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_1__6_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_1__7_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_1__8_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_1__9_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_1__10_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_1__11_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_1__12_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_1__13_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_2__0_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_2__1_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_2__2_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_2__3_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_2__4_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_2__5_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_2__6_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_2__7_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_2__8_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_2__9_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_2__10_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_2__11_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_2__12_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_2__13_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_3__0_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_3__1_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_3__2_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_3__3_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_3__4_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_3__5_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_3__6_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_3__7_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_3__8_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_3__9_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_3__10_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_3__11_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_3__12_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_3__13_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_4__0_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_4__1_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_4__2_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_4__3_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_4__4_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_4__5_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_4__6_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_4__7_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_4__8_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_4__9_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_4__10_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_4__11_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_4__12_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_4__13_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_5__0_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_5__1_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_5__2_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_5__3_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_5__4_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_5__5_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_5__6_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_5__7_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_5__8_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_5__9_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_5__10_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_5__11_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_5__12_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_5__13_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_6__0_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_6__1_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_6__2_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_6__3_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_6__4_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_6__5_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_6__6_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_6__7_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_6__8_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_6__9_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_6__10_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_6__11_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_6__12_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_6__13_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_7__0_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_7__1_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_7__2_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_7__3_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_7__4_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_7__5_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_7__6_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_7__7_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_7__8_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_7__9_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_7__10_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_7__11_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_7__12_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_7__13_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_8__0_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_8__1_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_8__2_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_8__3_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_8__4_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_8__5_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_8__6_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_8__7_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_8__8_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_8__9_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_8__10_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_8__11_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_8__12_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_8__13_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_9__0_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_9__1_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_9__2_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_9__3_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_9__4_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_9__5_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_9__6_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_9__7_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_9__8_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_9__9_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_9__10_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_9__11_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_9__12_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_9__13_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_10__0_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_10__1_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_10__2_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_10__3_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_10__4_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_10__5_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_10__6_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_10__7_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_10__8_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_10__9_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_10__10_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_10__11_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_10__12_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_10__13_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_11__0_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_11__1_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_11__2_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_11__3_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_11__4_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_11__5_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_11__6_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_11__7_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_11__8_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_11__9_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_11__10_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_11__11_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_11__12_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_11__13_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_12__0_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_12__1_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_12__2_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_12__3_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_12__4_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_12__5_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_12__6_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_12__7_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_12__8_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_12__9_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_12__10_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_12__11_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_12__12_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_12__13_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_13__0_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_13__1_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_13__2_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_13__3_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_13__4_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_13__5_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_13__6_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_13__7_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_13__8_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_13__9_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_13__10_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_13__11_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_13__12_,
         my_filter_adder_mult_7_multiplication_mult_21_ab_13__13_,
         my_filter_adder_mult_7_multiplication_mult_21_FS_1_n71,
         my_filter_adder_mult_7_multiplication_mult_21_FS_1_n70,
         my_filter_adder_mult_7_multiplication_mult_21_FS_1_n69,
         my_filter_adder_mult_7_multiplication_mult_21_FS_1_n68,
         my_filter_adder_mult_7_multiplication_mult_21_FS_1_n67,
         my_filter_adder_mult_7_multiplication_mult_21_FS_1_n66,
         my_filter_adder_mult_7_multiplication_mult_21_FS_1_n65,
         my_filter_adder_mult_7_multiplication_mult_21_FS_1_n64,
         my_filter_adder_mult_7_multiplication_mult_21_FS_1_n63,
         my_filter_adder_mult_7_multiplication_mult_21_FS_1_n62,
         my_filter_adder_mult_7_multiplication_mult_21_FS_1_n60,
         my_filter_adder_mult_7_multiplication_mult_21_FS_1_n59,
         my_filter_adder_mult_7_multiplication_mult_21_FS_1_n58,
         my_filter_adder_mult_7_multiplication_mult_21_FS_1_n57,
         my_filter_adder_mult_7_multiplication_mult_21_FS_1_n56,
         my_filter_adder_mult_7_multiplication_mult_21_FS_1_n55,
         my_filter_adder_mult_7_multiplication_mult_21_FS_1_n54,
         my_filter_adder_mult_7_multiplication_mult_21_FS_1_n53,
         my_filter_adder_mult_7_multiplication_mult_21_FS_1_n52,
         my_filter_adder_mult_7_multiplication_mult_21_FS_1_n51,
         my_filter_adder_mult_7_multiplication_mult_21_FS_1_n50,
         my_filter_adder_mult_7_multiplication_mult_21_FS_1_n49,
         my_filter_adder_mult_7_multiplication_mult_21_FS_1_n48,
         my_filter_adder_mult_7_multiplication_mult_21_FS_1_n47,
         my_filter_adder_mult_7_multiplication_mult_21_FS_1_n46,
         my_filter_adder_mult_7_multiplication_mult_21_FS_1_n45,
         my_filter_adder_mult_7_multiplication_mult_21_FS_1_n44,
         my_filter_adder_mult_7_multiplication_mult_21_FS_1_n43,
         my_filter_adder_mult_7_multiplication_mult_21_FS_1_n42,
         my_filter_adder_mult_7_multiplication_mult_21_FS_1_n41,
         my_filter_adder_mult_7_multiplication_mult_21_FS_1_n40,
         my_filter_adder_mult_7_multiplication_mult_21_FS_1_n39,
         my_filter_adder_mult_7_multiplication_mult_21_FS_1_n38,
         my_filter_adder_mult_7_multiplication_mult_21_FS_1_n37,
         my_filter_adder_mult_7_multiplication_mult_21_FS_1_n36,
         my_filter_adder_mult_7_multiplication_mult_21_FS_1_n35,
         my_filter_adder_mult_7_multiplication_mult_21_FS_1_n34,
         my_filter_adder_mult_7_multiplication_mult_21_FS_1_n33,
         my_filter_adder_mult_7_multiplication_mult_21_FS_1_n32,
         my_filter_adder_mult_7_multiplication_mult_21_FS_1_n31,
         my_filter_adder_mult_7_multiplication_mult_21_FS_1_n30,
         my_filter_adder_mult_7_multiplication_mult_21_FS_1_n29,
         my_filter_adder_mult_7_multiplication_mult_21_FS_1_n28,
         my_filter_adder_mult_7_multiplication_mult_21_FS_1_n27,
         my_filter_adder_mult_7_multiplication_mult_21_FS_1_n26,
         my_filter_adder_mult_7_multiplication_mult_21_FS_1_n25,
         my_filter_adder_mult_7_multiplication_mult_21_FS_1_n24,
         my_filter_adder_mult_7_multiplication_mult_21_FS_1_n23,
         my_filter_adder_mult_7_multiplication_mult_21_FS_1_n22,
         my_filter_adder_mult_7_multiplication_mult_21_FS_1_n21,
         my_filter_adder_mult_7_multiplication_mult_21_FS_1_n20,
         my_filter_adder_mult_7_multiplication_mult_21_FS_1_n19,
         my_filter_adder_mult_7_multiplication_mult_21_FS_1_n18,
         my_filter_adder_mult_7_multiplication_mult_21_FS_1_n17,
         my_filter_adder_mult_7_multiplication_mult_21_FS_1_n16,
         my_filter_adder_mult_7_multiplication_mult_21_FS_1_n15,
         my_filter_adder_mult_7_multiplication_mult_21_FS_1_n14,
         my_filter_adder_mult_7_multiplication_mult_21_FS_1_n13,
         my_filter_adder_mult_7_addition_add_19_n1,
         my_filter_adder_mult_8_multiplication_mult_21_n113,
         my_filter_adder_mult_8_multiplication_mult_21_n112,
         my_filter_adder_mult_8_multiplication_mult_21_n111,
         my_filter_adder_mult_8_multiplication_mult_21_n110,
         my_filter_adder_mult_8_multiplication_mult_21_n109,
         my_filter_adder_mult_8_multiplication_mult_21_n108,
         my_filter_adder_mult_8_multiplication_mult_21_n107,
         my_filter_adder_mult_8_multiplication_mult_21_n106,
         my_filter_adder_mult_8_multiplication_mult_21_n105,
         my_filter_adder_mult_8_multiplication_mult_21_n104,
         my_filter_adder_mult_8_multiplication_mult_21_n103,
         my_filter_adder_mult_8_multiplication_mult_21_n102,
         my_filter_adder_mult_8_multiplication_mult_21_n101,
         my_filter_adder_mult_8_multiplication_mult_21_n100,
         my_filter_adder_mult_8_multiplication_mult_21_n99,
         my_filter_adder_mult_8_multiplication_mult_21_n98,
         my_filter_adder_mult_8_multiplication_mult_21_n97,
         my_filter_adder_mult_8_multiplication_mult_21_n96,
         my_filter_adder_mult_8_multiplication_mult_21_n95,
         my_filter_adder_mult_8_multiplication_mult_21_n94,
         my_filter_adder_mult_8_multiplication_mult_21_n93,
         my_filter_adder_mult_8_multiplication_mult_21_n92,
         my_filter_adder_mult_8_multiplication_mult_21_n91,
         my_filter_adder_mult_8_multiplication_mult_21_n90,
         my_filter_adder_mult_8_multiplication_mult_21_n89,
         my_filter_adder_mult_8_multiplication_mult_21_n88,
         my_filter_adder_mult_8_multiplication_mult_21_n87,
         my_filter_adder_mult_8_multiplication_mult_21_n86,
         my_filter_adder_mult_8_multiplication_mult_21_n85,
         my_filter_adder_mult_8_multiplication_mult_21_n52,
         my_filter_adder_mult_8_multiplication_mult_21_n51,
         my_filter_adder_mult_8_multiplication_mult_21_n50,
         my_filter_adder_mult_8_multiplication_mult_21_n49,
         my_filter_adder_mult_8_multiplication_mult_21_n48,
         my_filter_adder_mult_8_multiplication_mult_21_n47,
         my_filter_adder_mult_8_multiplication_mult_21_n46,
         my_filter_adder_mult_8_multiplication_mult_21_n45,
         my_filter_adder_mult_8_multiplication_mult_21_n44,
         my_filter_adder_mult_8_multiplication_mult_21_n43,
         my_filter_adder_mult_8_multiplication_mult_21_n42,
         my_filter_adder_mult_8_multiplication_mult_21_n41,
         my_filter_adder_mult_8_multiplication_mult_21_n40,
         my_filter_adder_mult_8_multiplication_mult_21_n39,
         my_filter_adder_mult_8_multiplication_mult_21_n38,
         my_filter_adder_mult_8_multiplication_mult_21_n37,
         my_filter_adder_mult_8_multiplication_mult_21_n36,
         my_filter_adder_mult_8_multiplication_mult_21_n35,
         my_filter_adder_mult_8_multiplication_mult_21_n34,
         my_filter_adder_mult_8_multiplication_mult_21_n33,
         my_filter_adder_mult_8_multiplication_mult_21_n32,
         my_filter_adder_mult_8_multiplication_mult_21_n31,
         my_filter_adder_mult_8_multiplication_mult_21_n30,
         my_filter_adder_mult_8_multiplication_mult_21_n29,
         my_filter_adder_mult_8_multiplication_mult_21_n28,
         my_filter_adder_mult_8_multiplication_mult_21_n27,
         my_filter_adder_mult_8_multiplication_mult_21_n26,
         my_filter_adder_mult_8_multiplication_mult_21_n25,
         my_filter_adder_mult_8_multiplication_mult_21_n24,
         my_filter_adder_mult_8_multiplication_mult_21_n23,
         my_filter_adder_mult_8_multiplication_mult_21_n22,
         my_filter_adder_mult_8_multiplication_mult_21_n21,
         my_filter_adder_mult_8_multiplication_mult_21_n20,
         my_filter_adder_mult_8_multiplication_mult_21_n19,
         my_filter_adder_mult_8_multiplication_mult_21_n18,
         my_filter_adder_mult_8_multiplication_mult_21_n17,
         my_filter_adder_mult_8_multiplication_mult_21_n16,
         my_filter_adder_mult_8_multiplication_mult_21_n15,
         my_filter_adder_mult_8_multiplication_mult_21_n14,
         my_filter_adder_mult_8_multiplication_mult_21_n13,
         my_filter_adder_mult_8_multiplication_mult_21_n12,
         my_filter_adder_mult_8_multiplication_mult_21_n11,
         my_filter_adder_mult_8_multiplication_mult_21_n10,
         my_filter_adder_mult_8_multiplication_mult_21_n9,
         my_filter_adder_mult_8_multiplication_mult_21_n8,
         my_filter_adder_mult_8_multiplication_mult_21_n7,
         my_filter_adder_mult_8_multiplication_mult_21_n6,
         my_filter_adder_mult_8_multiplication_mult_21_n5,
         my_filter_adder_mult_8_multiplication_mult_21_n4,
         my_filter_adder_mult_8_multiplication_mult_21_n3,
         my_filter_adder_mult_8_multiplication_mult_21_A2_12_,
         my_filter_adder_mult_8_multiplication_mult_21_A1_0_,
         my_filter_adder_mult_8_multiplication_mult_21_A1_1_,
         my_filter_adder_mult_8_multiplication_mult_21_A1_2_,
         my_filter_adder_mult_8_multiplication_mult_21_A1_3_,
         my_filter_adder_mult_8_multiplication_mult_21_A1_4_,
         my_filter_adder_mult_8_multiplication_mult_21_A1_5_,
         my_filter_adder_mult_8_multiplication_mult_21_A1_6_,
         my_filter_adder_mult_8_multiplication_mult_21_A1_7_,
         my_filter_adder_mult_8_multiplication_mult_21_A1_8_,
         my_filter_adder_mult_8_multiplication_mult_21_A1_9_,
         my_filter_adder_mult_8_multiplication_mult_21_A1_10_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_2__1_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_2__2_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_2__3_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_2__4_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_2__5_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_2__6_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_2__7_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_2__8_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_2__9_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_2__10_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_2__11_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_2__12_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_3__1_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_3__2_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_3__3_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_3__4_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_3__5_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_3__6_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_3__7_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_3__8_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_3__9_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_3__10_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_3__11_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_3__12_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_4__1_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_4__2_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_4__3_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_4__4_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_4__5_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_4__6_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_4__7_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_4__8_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_4__9_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_4__10_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_4__11_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_4__12_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_5__1_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_5__2_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_5__3_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_5__4_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_5__5_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_5__6_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_5__7_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_5__8_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_5__9_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_5__10_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_5__11_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_5__12_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_6__1_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_6__2_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_6__3_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_6__4_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_6__5_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_6__6_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_6__7_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_6__8_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_6__9_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_6__10_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_6__11_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_6__12_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_7__1_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_7__2_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_7__3_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_7__4_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_7__5_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_7__6_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_7__7_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_7__8_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_7__9_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_7__10_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_7__11_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_7__12_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_8__1_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_8__2_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_8__3_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_8__4_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_8__5_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_8__6_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_8__7_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_8__8_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_8__9_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_8__10_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_8__11_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_8__12_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_9__1_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_9__2_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_9__3_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_9__4_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_9__5_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_9__6_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_9__7_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_9__8_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_9__9_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_9__10_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_9__11_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_9__12_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_10__1_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_10__2_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_10__3_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_10__4_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_10__5_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_10__6_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_10__7_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_10__8_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_10__9_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_10__10_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_10__11_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_10__12_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_11__1_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_11__2_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_11__3_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_11__4_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_11__5_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_11__6_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_11__7_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_11__8_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_11__9_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_11__10_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_11__11_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_11__12_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_12__1_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_12__2_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_12__3_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_12__4_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_12__5_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_12__6_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_12__7_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_12__8_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_12__9_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_12__10_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_12__11_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_12__12_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_13__0_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_13__1_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_13__2_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_13__3_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_13__4_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_13__5_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_13__6_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_13__7_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_13__8_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_13__9_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_13__10_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_13__11_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_13__12_,
         my_filter_adder_mult_8_multiplication_mult_21_SUMB_13__13_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_1__0_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_2__0_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_2__1_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_2__2_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_2__3_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_2__4_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_2__5_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_2__6_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_2__7_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_2__8_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_2__9_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_2__10_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_2__11_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_2__12_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_3__0_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_3__1_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_3__2_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_3__3_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_3__4_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_3__5_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_3__6_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_3__7_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_3__8_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_3__9_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_3__10_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_3__11_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_3__12_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_4__0_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_4__1_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_4__2_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_4__3_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_4__4_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_4__5_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_4__6_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_4__7_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_4__8_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_4__9_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_4__10_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_4__11_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_4__12_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_5__0_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_5__1_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_5__2_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_5__3_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_5__4_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_5__5_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_5__6_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_5__7_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_5__8_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_5__9_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_5__10_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_5__11_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_5__12_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_6__0_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_6__1_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_6__2_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_6__3_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_6__4_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_6__5_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_6__6_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_6__7_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_6__8_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_6__9_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_6__10_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_6__11_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_6__12_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_7__0_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_7__1_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_7__2_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_7__3_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_7__4_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_7__5_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_7__6_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_7__7_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_7__8_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_7__9_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_7__10_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_7__11_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_7__12_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_8__0_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_8__1_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_8__2_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_8__3_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_8__4_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_8__5_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_8__6_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_8__7_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_8__8_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_8__9_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_8__10_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_8__11_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_8__12_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_9__0_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_9__1_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_9__2_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_9__3_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_9__4_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_9__5_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_9__6_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_9__7_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_9__8_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_9__9_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_9__10_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_9__11_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_9__12_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_10__0_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_10__1_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_10__2_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_10__3_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_10__4_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_10__5_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_10__6_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_10__7_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_10__8_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_10__9_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_10__10_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_10__11_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_10__12_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_11__0_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_11__1_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_11__2_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_11__3_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_11__4_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_11__5_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_11__6_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_11__7_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_11__8_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_11__9_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_11__10_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_11__11_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_11__12_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_12__0_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_12__1_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_12__2_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_12__3_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_12__4_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_12__5_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_12__6_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_12__7_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_12__8_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_12__9_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_12__10_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_12__11_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_12__12_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_13__0_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_13__1_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_13__2_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_13__3_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_13__4_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_13__5_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_13__6_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_13__7_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_13__8_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_13__9_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_13__10_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_13__11_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_13__12_,
         my_filter_adder_mult_8_multiplication_mult_21_CARRYB_13__13_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_0__2_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_0__3_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_0__4_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_0__5_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_0__6_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_0__7_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_0__8_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_0__9_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_0__10_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_0__11_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_0__12_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_0__13_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_1__1_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_1__2_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_1__3_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_1__4_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_1__5_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_1__6_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_1__7_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_1__8_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_1__9_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_1__10_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_1__11_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_1__12_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_1__13_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_2__0_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_2__1_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_2__2_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_2__3_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_2__4_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_2__5_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_2__6_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_2__7_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_2__8_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_2__9_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_2__10_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_2__11_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_2__12_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_2__13_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_3__0_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_3__1_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_3__2_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_3__3_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_3__4_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_3__5_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_3__6_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_3__7_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_3__8_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_3__9_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_3__10_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_3__11_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_3__12_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_3__13_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_4__0_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_4__1_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_4__2_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_4__3_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_4__4_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_4__5_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_4__6_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_4__7_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_4__8_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_4__9_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_4__10_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_4__11_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_4__12_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_4__13_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_5__0_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_5__1_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_5__2_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_5__3_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_5__4_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_5__5_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_5__6_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_5__7_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_5__8_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_5__9_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_5__10_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_5__11_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_5__12_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_5__13_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_6__0_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_6__1_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_6__2_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_6__3_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_6__4_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_6__5_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_6__6_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_6__7_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_6__8_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_6__9_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_6__10_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_6__11_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_6__12_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_6__13_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_7__0_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_7__1_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_7__2_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_7__3_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_7__4_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_7__5_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_7__6_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_7__7_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_7__8_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_7__9_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_7__10_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_7__11_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_7__12_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_7__13_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_8__0_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_8__1_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_8__2_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_8__3_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_8__4_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_8__5_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_8__6_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_8__7_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_8__8_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_8__9_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_8__10_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_8__11_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_8__12_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_8__13_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_9__0_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_9__1_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_9__2_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_9__3_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_9__4_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_9__5_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_9__6_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_9__7_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_9__8_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_9__9_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_9__10_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_9__11_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_9__12_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_9__13_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_10__0_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_10__1_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_10__2_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_10__3_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_10__4_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_10__5_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_10__6_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_10__7_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_10__8_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_10__9_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_10__10_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_10__11_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_10__12_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_10__13_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_11__0_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_11__1_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_11__2_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_11__3_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_11__4_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_11__5_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_11__6_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_11__7_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_11__8_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_11__9_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_11__10_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_11__11_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_11__12_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_11__13_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_12__0_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_12__1_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_12__2_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_12__3_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_12__4_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_12__5_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_12__6_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_12__7_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_12__8_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_12__9_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_12__10_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_12__11_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_12__12_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_12__13_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_13__0_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_13__1_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_13__2_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_13__3_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_13__4_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_13__5_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_13__6_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_13__7_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_13__8_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_13__9_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_13__10_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_13__11_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_13__12_,
         my_filter_adder_mult_8_multiplication_mult_21_ab_13__13_,
         my_filter_adder_mult_8_multiplication_mult_21_FS_1_n71,
         my_filter_adder_mult_8_multiplication_mult_21_FS_1_n70,
         my_filter_adder_mult_8_multiplication_mult_21_FS_1_n69,
         my_filter_adder_mult_8_multiplication_mult_21_FS_1_n68,
         my_filter_adder_mult_8_multiplication_mult_21_FS_1_n67,
         my_filter_adder_mult_8_multiplication_mult_21_FS_1_n66,
         my_filter_adder_mult_8_multiplication_mult_21_FS_1_n65,
         my_filter_adder_mult_8_multiplication_mult_21_FS_1_n64,
         my_filter_adder_mult_8_multiplication_mult_21_FS_1_n63,
         my_filter_adder_mult_8_multiplication_mult_21_FS_1_n62,
         my_filter_adder_mult_8_multiplication_mult_21_FS_1_n60,
         my_filter_adder_mult_8_multiplication_mult_21_FS_1_n59,
         my_filter_adder_mult_8_multiplication_mult_21_FS_1_n58,
         my_filter_adder_mult_8_multiplication_mult_21_FS_1_n57,
         my_filter_adder_mult_8_multiplication_mult_21_FS_1_n56,
         my_filter_adder_mult_8_multiplication_mult_21_FS_1_n55,
         my_filter_adder_mult_8_multiplication_mult_21_FS_1_n54,
         my_filter_adder_mult_8_multiplication_mult_21_FS_1_n53,
         my_filter_adder_mult_8_multiplication_mult_21_FS_1_n52,
         my_filter_adder_mult_8_multiplication_mult_21_FS_1_n51,
         my_filter_adder_mult_8_multiplication_mult_21_FS_1_n50,
         my_filter_adder_mult_8_multiplication_mult_21_FS_1_n49,
         my_filter_adder_mult_8_multiplication_mult_21_FS_1_n48,
         my_filter_adder_mult_8_multiplication_mult_21_FS_1_n47,
         my_filter_adder_mult_8_multiplication_mult_21_FS_1_n46,
         my_filter_adder_mult_8_multiplication_mult_21_FS_1_n45,
         my_filter_adder_mult_8_multiplication_mult_21_FS_1_n44,
         my_filter_adder_mult_8_multiplication_mult_21_FS_1_n43,
         my_filter_adder_mult_8_multiplication_mult_21_FS_1_n42,
         my_filter_adder_mult_8_multiplication_mult_21_FS_1_n41,
         my_filter_adder_mult_8_multiplication_mult_21_FS_1_n40,
         my_filter_adder_mult_8_multiplication_mult_21_FS_1_n39,
         my_filter_adder_mult_8_multiplication_mult_21_FS_1_n38,
         my_filter_adder_mult_8_multiplication_mult_21_FS_1_n37,
         my_filter_adder_mult_8_multiplication_mult_21_FS_1_n36,
         my_filter_adder_mult_8_multiplication_mult_21_FS_1_n35,
         my_filter_adder_mult_8_multiplication_mult_21_FS_1_n34,
         my_filter_adder_mult_8_multiplication_mult_21_FS_1_n33,
         my_filter_adder_mult_8_multiplication_mult_21_FS_1_n32,
         my_filter_adder_mult_8_multiplication_mult_21_FS_1_n31,
         my_filter_adder_mult_8_multiplication_mult_21_FS_1_n30,
         my_filter_adder_mult_8_multiplication_mult_21_FS_1_n29,
         my_filter_adder_mult_8_multiplication_mult_21_FS_1_n28,
         my_filter_adder_mult_8_multiplication_mult_21_FS_1_n27,
         my_filter_adder_mult_8_multiplication_mult_21_FS_1_n26,
         my_filter_adder_mult_8_multiplication_mult_21_FS_1_n25,
         my_filter_adder_mult_8_multiplication_mult_21_FS_1_n24,
         my_filter_adder_mult_8_multiplication_mult_21_FS_1_n23,
         my_filter_adder_mult_8_multiplication_mult_21_FS_1_n22,
         my_filter_adder_mult_8_multiplication_mult_21_FS_1_n21,
         my_filter_adder_mult_8_multiplication_mult_21_FS_1_n20,
         my_filter_adder_mult_8_multiplication_mult_21_FS_1_n19,
         my_filter_adder_mult_8_multiplication_mult_21_FS_1_n18,
         my_filter_adder_mult_8_multiplication_mult_21_FS_1_n17,
         my_filter_adder_mult_8_multiplication_mult_21_FS_1_n16,
         my_filter_adder_mult_8_multiplication_mult_21_FS_1_n15,
         my_filter_adder_mult_8_multiplication_mult_21_FS_1_n14,
         my_filter_adder_mult_8_multiplication_mult_21_FS_1_n13,
         my_filter_adder_mult_8_addition_add_19_n1,
         my_filter_adder_mult_9_multiplication_mult_21_n113,
         my_filter_adder_mult_9_multiplication_mult_21_n112,
         my_filter_adder_mult_9_multiplication_mult_21_n111,
         my_filter_adder_mult_9_multiplication_mult_21_n110,
         my_filter_adder_mult_9_multiplication_mult_21_n109,
         my_filter_adder_mult_9_multiplication_mult_21_n108,
         my_filter_adder_mult_9_multiplication_mult_21_n107,
         my_filter_adder_mult_9_multiplication_mult_21_n106,
         my_filter_adder_mult_9_multiplication_mult_21_n105,
         my_filter_adder_mult_9_multiplication_mult_21_n104,
         my_filter_adder_mult_9_multiplication_mult_21_n103,
         my_filter_adder_mult_9_multiplication_mult_21_n102,
         my_filter_adder_mult_9_multiplication_mult_21_n101,
         my_filter_adder_mult_9_multiplication_mult_21_n100,
         my_filter_adder_mult_9_multiplication_mult_21_n99,
         my_filter_adder_mult_9_multiplication_mult_21_n98,
         my_filter_adder_mult_9_multiplication_mult_21_n97,
         my_filter_adder_mult_9_multiplication_mult_21_n96,
         my_filter_adder_mult_9_multiplication_mult_21_n95,
         my_filter_adder_mult_9_multiplication_mult_21_n94,
         my_filter_adder_mult_9_multiplication_mult_21_n93,
         my_filter_adder_mult_9_multiplication_mult_21_n92,
         my_filter_adder_mult_9_multiplication_mult_21_n91,
         my_filter_adder_mult_9_multiplication_mult_21_n90,
         my_filter_adder_mult_9_multiplication_mult_21_n89,
         my_filter_adder_mult_9_multiplication_mult_21_n88,
         my_filter_adder_mult_9_multiplication_mult_21_n87,
         my_filter_adder_mult_9_multiplication_mult_21_n86,
         my_filter_adder_mult_9_multiplication_mult_21_n85,
         my_filter_adder_mult_9_multiplication_mult_21_n52,
         my_filter_adder_mult_9_multiplication_mult_21_n51,
         my_filter_adder_mult_9_multiplication_mult_21_n50,
         my_filter_adder_mult_9_multiplication_mult_21_n49,
         my_filter_adder_mult_9_multiplication_mult_21_n48,
         my_filter_adder_mult_9_multiplication_mult_21_n47,
         my_filter_adder_mult_9_multiplication_mult_21_n46,
         my_filter_adder_mult_9_multiplication_mult_21_n45,
         my_filter_adder_mult_9_multiplication_mult_21_n44,
         my_filter_adder_mult_9_multiplication_mult_21_n43,
         my_filter_adder_mult_9_multiplication_mult_21_n42,
         my_filter_adder_mult_9_multiplication_mult_21_n41,
         my_filter_adder_mult_9_multiplication_mult_21_n40,
         my_filter_adder_mult_9_multiplication_mult_21_n39,
         my_filter_adder_mult_9_multiplication_mult_21_n38,
         my_filter_adder_mult_9_multiplication_mult_21_n37,
         my_filter_adder_mult_9_multiplication_mult_21_n36,
         my_filter_adder_mult_9_multiplication_mult_21_n35,
         my_filter_adder_mult_9_multiplication_mult_21_n34,
         my_filter_adder_mult_9_multiplication_mult_21_n33,
         my_filter_adder_mult_9_multiplication_mult_21_n32,
         my_filter_adder_mult_9_multiplication_mult_21_n31,
         my_filter_adder_mult_9_multiplication_mult_21_n30,
         my_filter_adder_mult_9_multiplication_mult_21_n29,
         my_filter_adder_mult_9_multiplication_mult_21_n28,
         my_filter_adder_mult_9_multiplication_mult_21_n27,
         my_filter_adder_mult_9_multiplication_mult_21_n26,
         my_filter_adder_mult_9_multiplication_mult_21_n25,
         my_filter_adder_mult_9_multiplication_mult_21_n24,
         my_filter_adder_mult_9_multiplication_mult_21_n23,
         my_filter_adder_mult_9_multiplication_mult_21_n22,
         my_filter_adder_mult_9_multiplication_mult_21_n21,
         my_filter_adder_mult_9_multiplication_mult_21_n20,
         my_filter_adder_mult_9_multiplication_mult_21_n19,
         my_filter_adder_mult_9_multiplication_mult_21_n18,
         my_filter_adder_mult_9_multiplication_mult_21_n17,
         my_filter_adder_mult_9_multiplication_mult_21_n16,
         my_filter_adder_mult_9_multiplication_mult_21_n15,
         my_filter_adder_mult_9_multiplication_mult_21_n14,
         my_filter_adder_mult_9_multiplication_mult_21_n13,
         my_filter_adder_mult_9_multiplication_mult_21_n12,
         my_filter_adder_mult_9_multiplication_mult_21_n11,
         my_filter_adder_mult_9_multiplication_mult_21_n10,
         my_filter_adder_mult_9_multiplication_mult_21_n9,
         my_filter_adder_mult_9_multiplication_mult_21_n8,
         my_filter_adder_mult_9_multiplication_mult_21_n7,
         my_filter_adder_mult_9_multiplication_mult_21_n6,
         my_filter_adder_mult_9_multiplication_mult_21_n5,
         my_filter_adder_mult_9_multiplication_mult_21_n4,
         my_filter_adder_mult_9_multiplication_mult_21_n3,
         my_filter_adder_mult_9_multiplication_mult_21_A2_12_,
         my_filter_adder_mult_9_multiplication_mult_21_A1_0_,
         my_filter_adder_mult_9_multiplication_mult_21_A1_1_,
         my_filter_adder_mult_9_multiplication_mult_21_A1_2_,
         my_filter_adder_mult_9_multiplication_mult_21_A1_3_,
         my_filter_adder_mult_9_multiplication_mult_21_A1_4_,
         my_filter_adder_mult_9_multiplication_mult_21_A1_5_,
         my_filter_adder_mult_9_multiplication_mult_21_A1_6_,
         my_filter_adder_mult_9_multiplication_mult_21_A1_7_,
         my_filter_adder_mult_9_multiplication_mult_21_A1_8_,
         my_filter_adder_mult_9_multiplication_mult_21_A1_9_,
         my_filter_adder_mult_9_multiplication_mult_21_A1_10_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_2__1_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_2__2_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_2__3_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_2__4_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_2__5_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_2__6_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_2__7_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_2__8_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_2__9_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_2__10_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_2__11_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_2__12_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_3__1_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_3__2_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_3__3_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_3__4_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_3__5_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_3__6_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_3__7_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_3__8_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_3__9_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_3__10_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_3__11_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_3__12_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_4__1_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_4__2_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_4__3_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_4__4_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_4__5_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_4__6_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_4__7_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_4__8_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_4__9_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_4__10_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_4__11_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_4__12_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_5__1_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_5__2_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_5__3_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_5__4_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_5__5_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_5__6_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_5__7_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_5__8_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_5__9_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_5__10_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_5__11_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_5__12_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_6__1_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_6__2_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_6__3_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_6__4_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_6__5_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_6__6_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_6__7_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_6__8_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_6__9_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_6__10_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_6__11_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_6__12_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_7__1_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_7__2_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_7__3_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_7__4_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_7__5_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_7__6_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_7__7_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_7__8_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_7__9_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_7__10_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_7__11_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_7__12_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_8__1_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_8__2_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_8__3_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_8__4_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_8__5_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_8__6_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_8__7_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_8__8_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_8__9_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_8__10_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_8__11_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_8__12_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_9__1_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_9__2_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_9__3_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_9__4_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_9__5_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_9__6_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_9__7_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_9__8_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_9__9_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_9__10_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_9__11_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_9__12_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_10__1_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_10__2_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_10__3_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_10__4_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_10__5_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_10__6_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_10__7_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_10__8_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_10__9_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_10__10_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_10__11_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_10__12_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_11__1_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_11__2_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_11__3_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_11__4_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_11__5_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_11__6_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_11__7_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_11__8_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_11__9_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_11__10_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_11__11_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_11__12_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_12__1_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_12__2_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_12__3_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_12__4_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_12__5_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_12__6_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_12__7_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_12__8_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_12__9_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_12__10_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_12__11_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_12__12_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_13__0_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_13__1_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_13__2_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_13__3_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_13__4_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_13__5_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_13__6_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_13__7_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_13__8_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_13__9_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_13__10_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_13__11_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_13__12_,
         my_filter_adder_mult_9_multiplication_mult_21_SUMB_13__13_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_1__0_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_2__0_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_2__1_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_2__2_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_2__3_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_2__4_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_2__5_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_2__6_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_2__7_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_2__8_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_2__9_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_2__10_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_2__11_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_2__12_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_3__0_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_3__1_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_3__2_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_3__3_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_3__4_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_3__5_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_3__6_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_3__7_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_3__8_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_3__9_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_3__10_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_3__11_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_3__12_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_4__0_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_4__1_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_4__2_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_4__3_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_4__4_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_4__5_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_4__6_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_4__7_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_4__8_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_4__9_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_4__10_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_4__11_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_4__12_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_5__0_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_5__1_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_5__2_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_5__3_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_5__4_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_5__5_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_5__6_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_5__7_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_5__8_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_5__9_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_5__10_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_5__11_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_5__12_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_6__0_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_6__1_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_6__2_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_6__3_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_6__4_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_6__5_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_6__6_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_6__7_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_6__8_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_6__9_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_6__10_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_6__11_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_6__12_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_7__0_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_7__1_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_7__2_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_7__3_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_7__4_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_7__5_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_7__6_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_7__7_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_7__8_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_7__9_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_7__10_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_7__11_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_7__12_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_8__0_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_8__1_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_8__2_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_8__3_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_8__4_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_8__5_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_8__6_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_8__7_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_8__8_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_8__9_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_8__10_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_8__11_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_8__12_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_9__0_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_9__1_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_9__2_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_9__3_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_9__4_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_9__5_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_9__6_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_9__7_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_9__8_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_9__9_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_9__10_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_9__11_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_9__12_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_10__0_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_10__1_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_10__2_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_10__3_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_10__4_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_10__5_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_10__6_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_10__7_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_10__8_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_10__9_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_10__10_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_10__11_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_10__12_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_11__0_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_11__1_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_11__2_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_11__3_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_11__4_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_11__5_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_11__6_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_11__7_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_11__8_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_11__9_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_11__10_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_11__11_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_11__12_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_12__0_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_12__1_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_12__2_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_12__3_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_12__4_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_12__5_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_12__6_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_12__7_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_12__8_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_12__9_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_12__10_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_12__11_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_12__12_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_13__0_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_13__1_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_13__2_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_13__3_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_13__4_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_13__5_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_13__6_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_13__7_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_13__8_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_13__9_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_13__10_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_13__11_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_13__12_,
         my_filter_adder_mult_9_multiplication_mult_21_CARRYB_13__13_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_0__2_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_0__3_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_0__4_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_0__5_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_0__6_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_0__7_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_0__8_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_0__9_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_0__10_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_0__11_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_0__12_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_0__13_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_1__1_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_1__2_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_1__3_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_1__4_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_1__5_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_1__6_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_1__7_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_1__8_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_1__9_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_1__10_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_1__11_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_1__12_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_1__13_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_2__0_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_2__1_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_2__2_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_2__3_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_2__4_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_2__5_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_2__6_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_2__7_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_2__8_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_2__9_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_2__10_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_2__11_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_2__12_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_2__13_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_3__0_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_3__1_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_3__2_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_3__3_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_3__4_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_3__5_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_3__6_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_3__7_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_3__8_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_3__9_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_3__10_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_3__11_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_3__12_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_3__13_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_4__0_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_4__1_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_4__2_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_4__3_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_4__4_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_4__5_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_4__6_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_4__7_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_4__8_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_4__9_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_4__10_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_4__11_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_4__12_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_4__13_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_5__0_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_5__1_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_5__2_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_5__3_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_5__4_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_5__5_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_5__6_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_5__7_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_5__8_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_5__9_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_5__10_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_5__11_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_5__12_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_5__13_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_6__0_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_6__1_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_6__2_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_6__3_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_6__4_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_6__5_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_6__6_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_6__7_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_6__8_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_6__9_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_6__10_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_6__11_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_6__12_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_6__13_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_7__0_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_7__1_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_7__2_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_7__3_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_7__4_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_7__5_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_7__6_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_7__7_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_7__8_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_7__9_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_7__10_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_7__11_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_7__12_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_7__13_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_8__0_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_8__1_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_8__2_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_8__3_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_8__4_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_8__5_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_8__6_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_8__7_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_8__8_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_8__9_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_8__10_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_8__11_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_8__12_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_8__13_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_9__0_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_9__1_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_9__2_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_9__3_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_9__4_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_9__5_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_9__6_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_9__7_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_9__8_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_9__9_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_9__10_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_9__11_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_9__12_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_9__13_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_10__0_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_10__1_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_10__2_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_10__3_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_10__4_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_10__5_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_10__6_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_10__7_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_10__8_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_10__9_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_10__10_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_10__11_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_10__12_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_10__13_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_11__0_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_11__1_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_11__2_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_11__3_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_11__4_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_11__5_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_11__6_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_11__7_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_11__8_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_11__9_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_11__10_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_11__11_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_11__12_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_11__13_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_12__0_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_12__1_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_12__2_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_12__3_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_12__4_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_12__5_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_12__6_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_12__7_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_12__8_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_12__9_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_12__10_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_12__11_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_12__12_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_12__13_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_13__0_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_13__1_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_13__2_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_13__3_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_13__4_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_13__5_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_13__6_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_13__7_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_13__8_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_13__9_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_13__10_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_13__11_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_13__12_,
         my_filter_adder_mult_9_multiplication_mult_21_ab_13__13_,
         my_filter_adder_mult_9_multiplication_mult_21_FS_1_n71,
         my_filter_adder_mult_9_multiplication_mult_21_FS_1_n70,
         my_filter_adder_mult_9_multiplication_mult_21_FS_1_n69,
         my_filter_adder_mult_9_multiplication_mult_21_FS_1_n68,
         my_filter_adder_mult_9_multiplication_mult_21_FS_1_n67,
         my_filter_adder_mult_9_multiplication_mult_21_FS_1_n66,
         my_filter_adder_mult_9_multiplication_mult_21_FS_1_n65,
         my_filter_adder_mult_9_multiplication_mult_21_FS_1_n64,
         my_filter_adder_mult_9_multiplication_mult_21_FS_1_n63,
         my_filter_adder_mult_9_multiplication_mult_21_FS_1_n62,
         my_filter_adder_mult_9_multiplication_mult_21_FS_1_n60,
         my_filter_adder_mult_9_multiplication_mult_21_FS_1_n59,
         my_filter_adder_mult_9_multiplication_mult_21_FS_1_n58,
         my_filter_adder_mult_9_multiplication_mult_21_FS_1_n57,
         my_filter_adder_mult_9_multiplication_mult_21_FS_1_n56,
         my_filter_adder_mult_9_multiplication_mult_21_FS_1_n55,
         my_filter_adder_mult_9_multiplication_mult_21_FS_1_n54,
         my_filter_adder_mult_9_multiplication_mult_21_FS_1_n53,
         my_filter_adder_mult_9_multiplication_mult_21_FS_1_n52,
         my_filter_adder_mult_9_multiplication_mult_21_FS_1_n51,
         my_filter_adder_mult_9_multiplication_mult_21_FS_1_n50,
         my_filter_adder_mult_9_multiplication_mult_21_FS_1_n49,
         my_filter_adder_mult_9_multiplication_mult_21_FS_1_n48,
         my_filter_adder_mult_9_multiplication_mult_21_FS_1_n47,
         my_filter_adder_mult_9_multiplication_mult_21_FS_1_n46,
         my_filter_adder_mult_9_multiplication_mult_21_FS_1_n45,
         my_filter_adder_mult_9_multiplication_mult_21_FS_1_n44,
         my_filter_adder_mult_9_multiplication_mult_21_FS_1_n43,
         my_filter_adder_mult_9_multiplication_mult_21_FS_1_n42,
         my_filter_adder_mult_9_multiplication_mult_21_FS_1_n41,
         my_filter_adder_mult_9_multiplication_mult_21_FS_1_n40,
         my_filter_adder_mult_9_multiplication_mult_21_FS_1_n39,
         my_filter_adder_mult_9_multiplication_mult_21_FS_1_n38,
         my_filter_adder_mult_9_multiplication_mult_21_FS_1_n37,
         my_filter_adder_mult_9_multiplication_mult_21_FS_1_n36,
         my_filter_adder_mult_9_multiplication_mult_21_FS_1_n35,
         my_filter_adder_mult_9_multiplication_mult_21_FS_1_n34,
         my_filter_adder_mult_9_multiplication_mult_21_FS_1_n33,
         my_filter_adder_mult_9_multiplication_mult_21_FS_1_n32,
         my_filter_adder_mult_9_multiplication_mult_21_FS_1_n31,
         my_filter_adder_mult_9_multiplication_mult_21_FS_1_n30,
         my_filter_adder_mult_9_multiplication_mult_21_FS_1_n29,
         my_filter_adder_mult_9_multiplication_mult_21_FS_1_n28,
         my_filter_adder_mult_9_multiplication_mult_21_FS_1_n27,
         my_filter_adder_mult_9_multiplication_mult_21_FS_1_n26,
         my_filter_adder_mult_9_multiplication_mult_21_FS_1_n25,
         my_filter_adder_mult_9_multiplication_mult_21_FS_1_n24,
         my_filter_adder_mult_9_multiplication_mult_21_FS_1_n23,
         my_filter_adder_mult_9_multiplication_mult_21_FS_1_n22,
         my_filter_adder_mult_9_multiplication_mult_21_FS_1_n21,
         my_filter_adder_mult_9_multiplication_mult_21_FS_1_n20,
         my_filter_adder_mult_9_multiplication_mult_21_FS_1_n19,
         my_filter_adder_mult_9_multiplication_mult_21_FS_1_n18,
         my_filter_adder_mult_9_multiplication_mult_21_FS_1_n17,
         my_filter_adder_mult_9_multiplication_mult_21_FS_1_n16,
         my_filter_adder_mult_9_multiplication_mult_21_FS_1_n15,
         my_filter_adder_mult_9_multiplication_mult_21_FS_1_n14,
         my_filter_adder_mult_9_multiplication_mult_21_FS_1_n13,
         my_filter_adder_mult_9_addition_add_19_n1;
  wire   [153:0] my_filter_data_sum;
  wire   [153:0] my_filter_q_reg_coeff;
  wire   [13:0] my_filter_adder_mult_0_res_mult;
  wire   [13:2] my_filter_adder_mult_0_addition_add_19_carry;
  wire   [13:0] my_filter_adder_mult_1_res_mult;
  wire   [13:2] my_filter_adder_mult_1_addition_add_19_carry;
  wire   [13:0] my_filter_adder_mult_2_res_mult;
  wire   [13:2] my_filter_adder_mult_2_addition_add_19_carry;
  wire   [13:0] my_filter_adder_mult_3_res_mult;
  wire   [13:2] my_filter_adder_mult_3_addition_add_19_carry;
  wire   [13:0] my_filter_adder_mult_4_res_mult;
  wire   [13:2] my_filter_adder_mult_4_addition_add_19_carry;
  wire   [13:0] my_filter_adder_mult_5_res_mult;
  wire   [13:2] my_filter_adder_mult_5_addition_add_19_carry;
  wire   [13:0] my_filter_adder_mult_6_res_mult;
  wire   [13:2] my_filter_adder_mult_6_addition_add_19_carry;
  wire   [13:0] my_filter_adder_mult_7_res_mult;
  wire   [13:2] my_filter_adder_mult_7_addition_add_19_carry;
  wire   [13:0] my_filter_adder_mult_8_res_mult;
  wire   [13:2] my_filter_adder_mult_8_addition_add_19_carry;
  wire   [13:0] my_filter_adder_mult_9_res_mult;
  wire   [13:2] my_filter_adder_mult_9_addition_add_19_carry;

  BUF_X1 my_filter_U1 ( .A(rst_n), .Z(my_filter_n2) );
  INV_X1 my_filter_reg_samples_U33 ( .A(vin), .ZN(my_filter_reg_samples_n45)
         );
  NAND2_X1 my_filter_reg_samples_U32 ( .A1(vin), .A2(din[13]), .ZN(
        my_filter_reg_samples_n3) );
  OAI21_X1 my_filter_reg_samples_U31 ( .B1(my_filter_reg_samples_n2), .B2(
        my_filter_reg_samples_n29), .A(my_filter_reg_samples_n3), .ZN(
        my_filter_reg_samples_n31) );
  NAND2_X1 my_filter_reg_samples_U30 ( .A1(din[12]), .A2(vin), .ZN(
        my_filter_reg_samples_n4) );
  OAI21_X1 my_filter_reg_samples_U29 ( .B1(my_filter_reg_samples_n2), .B2(
        my_filter_reg_samples_n28), .A(my_filter_reg_samples_n4), .ZN(
        my_filter_reg_samples_n32) );
  NAND2_X1 my_filter_reg_samples_U28 ( .A1(din[11]), .A2(vin), .ZN(
        my_filter_reg_samples_n5) );
  OAI21_X1 my_filter_reg_samples_U27 ( .B1(my_filter_reg_samples_n2), .B2(
        my_filter_reg_samples_n27), .A(my_filter_reg_samples_n5), .ZN(
        my_filter_reg_samples_n33) );
  NAND2_X1 my_filter_reg_samples_U26 ( .A1(din[10]), .A2(vin), .ZN(
        my_filter_reg_samples_n6) );
  OAI21_X1 my_filter_reg_samples_U25 ( .B1(my_filter_reg_samples_n2), .B2(
        my_filter_reg_samples_n26), .A(my_filter_reg_samples_n6), .ZN(
        my_filter_reg_samples_n34) );
  NAND2_X1 my_filter_reg_samples_U24 ( .A1(din[9]), .A2(vin), .ZN(
        my_filter_reg_samples_n7) );
  OAI21_X1 my_filter_reg_samples_U23 ( .B1(my_filter_reg_samples_n2), .B2(
        my_filter_reg_samples_n25), .A(my_filter_reg_samples_n7), .ZN(
        my_filter_reg_samples_n35) );
  NAND2_X1 my_filter_reg_samples_U22 ( .A1(din[8]), .A2(vin), .ZN(
        my_filter_reg_samples_n8) );
  OAI21_X1 my_filter_reg_samples_U21 ( .B1(my_filter_reg_samples_n2), .B2(
        my_filter_reg_samples_n24), .A(my_filter_reg_samples_n8), .ZN(
        my_filter_reg_samples_n36) );
  NAND2_X1 my_filter_reg_samples_U20 ( .A1(din[7]), .A2(vin), .ZN(
        my_filter_reg_samples_n9) );
  OAI21_X1 my_filter_reg_samples_U19 ( .B1(my_filter_reg_samples_n2), .B2(
        my_filter_reg_samples_n23), .A(my_filter_reg_samples_n9), .ZN(
        my_filter_reg_samples_n37) );
  NAND2_X1 my_filter_reg_samples_U18 ( .A1(din[6]), .A2(vin), .ZN(
        my_filter_reg_samples_n10) );
  OAI21_X1 my_filter_reg_samples_U17 ( .B1(my_filter_reg_samples_n2), .B2(
        my_filter_reg_samples_n22), .A(my_filter_reg_samples_n10), .ZN(
        my_filter_reg_samples_n38) );
  NAND2_X1 my_filter_reg_samples_U16 ( .A1(din[5]), .A2(vin), .ZN(
        my_filter_reg_samples_n11) );
  OAI21_X1 my_filter_reg_samples_U15 ( .B1(my_filter_reg_samples_n2), .B2(
        my_filter_reg_samples_n21), .A(my_filter_reg_samples_n11), .ZN(
        my_filter_reg_samples_n39) );
  NAND2_X1 my_filter_reg_samples_U14 ( .A1(din[4]), .A2(vin), .ZN(
        my_filter_reg_samples_n12) );
  OAI21_X1 my_filter_reg_samples_U13 ( .B1(my_filter_reg_samples_n2), .B2(
        my_filter_reg_samples_n20), .A(my_filter_reg_samples_n12), .ZN(
        my_filter_reg_samples_n40) );
  NAND2_X1 my_filter_reg_samples_U12 ( .A1(din[3]), .A2(vin), .ZN(
        my_filter_reg_samples_n13) );
  OAI21_X1 my_filter_reg_samples_U11 ( .B1(my_filter_reg_samples_n2), .B2(
        my_filter_reg_samples_n19), .A(my_filter_reg_samples_n13), .ZN(
        my_filter_reg_samples_n41) );
  NAND2_X1 my_filter_reg_samples_U10 ( .A1(din[2]), .A2(vin), .ZN(
        my_filter_reg_samples_n14) );
  OAI21_X1 my_filter_reg_samples_U9 ( .B1(my_filter_reg_samples_n2), .B2(
        my_filter_reg_samples_n18), .A(my_filter_reg_samples_n14), .ZN(
        my_filter_reg_samples_n42) );
  NAND2_X1 my_filter_reg_samples_U8 ( .A1(din[1]), .A2(vin), .ZN(
        my_filter_reg_samples_n15) );
  OAI21_X1 my_filter_reg_samples_U7 ( .B1(my_filter_reg_samples_n2), .B2(
        my_filter_reg_samples_n17), .A(my_filter_reg_samples_n15), .ZN(
        my_filter_reg_samples_n43) );
  NAND2_X1 my_filter_reg_samples_U6 ( .A1(din[0]), .A2(vin), .ZN(
        my_filter_reg_samples_n16) );
  OAI21_X1 my_filter_reg_samples_U5 ( .B1(my_filter_reg_samples_n2), .B2(
        my_filter_reg_samples_n30), .A(my_filter_reg_samples_n16), .ZN(
        my_filter_reg_samples_n44) );
  BUF_X1 my_filter_reg_samples_U4 ( .A(my_filter_n2), .Z(
        my_filter_reg_samples_n46) );
  NAND2_X1 my_filter_reg_samples_U3 ( .A1(my_filter_reg_samples_n46), .A2(
        my_filter_reg_samples_n45), .ZN(my_filter_reg_samples_n2) );
  DFFR_X1 my_filter_reg_samples_q_reg_0_ ( .D(my_filter_reg_samples_n44), .CK(
        clk), .RN(my_filter_reg_samples_n46), .Q(my_filter_q_reg_samp_0_), 
        .QN(my_filter_reg_samples_n30) );
  DFFR_X1 my_filter_reg_samples_q_reg_1_ ( .D(my_filter_reg_samples_n43), .CK(
        clk), .RN(my_filter_reg_samples_n46), .Q(my_filter_q_reg_samp_1_), 
        .QN(my_filter_reg_samples_n17) );
  DFFR_X1 my_filter_reg_samples_q_reg_2_ ( .D(my_filter_reg_samples_n42), .CK(
        clk), .RN(my_filter_reg_samples_n46), .Q(my_filter_q_reg_samp_2_), 
        .QN(my_filter_reg_samples_n18) );
  DFFR_X1 my_filter_reg_samples_q_reg_3_ ( .D(my_filter_reg_samples_n41), .CK(
        clk), .RN(my_filter_reg_samples_n46), .Q(my_filter_q_reg_samp_3_), 
        .QN(my_filter_reg_samples_n19) );
  DFFR_X1 my_filter_reg_samples_q_reg_4_ ( .D(my_filter_reg_samples_n40), .CK(
        clk), .RN(my_filter_reg_samples_n46), .Q(my_filter_q_reg_samp_4_), 
        .QN(my_filter_reg_samples_n20) );
  DFFR_X1 my_filter_reg_samples_q_reg_5_ ( .D(my_filter_reg_samples_n39), .CK(
        clk), .RN(my_filter_reg_samples_n46), .Q(my_filter_q_reg_samp_5_), 
        .QN(my_filter_reg_samples_n21) );
  DFFR_X1 my_filter_reg_samples_q_reg_6_ ( .D(my_filter_reg_samples_n38), .CK(
        clk), .RN(my_filter_reg_samples_n46), .Q(my_filter_q_reg_samp_6_), 
        .QN(my_filter_reg_samples_n22) );
  DFFR_X1 my_filter_reg_samples_q_reg_7_ ( .D(my_filter_reg_samples_n37), .CK(
        clk), .RN(my_filter_reg_samples_n46), .Q(my_filter_q_reg_samp_7_), 
        .QN(my_filter_reg_samples_n23) );
  DFFR_X1 my_filter_reg_samples_q_reg_8_ ( .D(my_filter_reg_samples_n36), .CK(
        clk), .RN(my_filter_reg_samples_n46), .Q(my_filter_q_reg_samp_8_), 
        .QN(my_filter_reg_samples_n24) );
  DFFR_X1 my_filter_reg_samples_q_reg_9_ ( .D(my_filter_reg_samples_n35), .CK(
        clk), .RN(my_filter_reg_samples_n46), .Q(my_filter_q_reg_samp_9_), 
        .QN(my_filter_reg_samples_n25) );
  DFFR_X1 my_filter_reg_samples_q_reg_10_ ( .D(my_filter_reg_samples_n34), 
        .CK(clk), .RN(my_filter_reg_samples_n46), .Q(my_filter_q_reg_samp_10_), 
        .QN(my_filter_reg_samples_n26) );
  DFFR_X1 my_filter_reg_samples_q_reg_11_ ( .D(my_filter_reg_samples_n33), 
        .CK(clk), .RN(my_filter_reg_samples_n46), .Q(my_filter_q_reg_samp_11_), 
        .QN(my_filter_reg_samples_n27) );
  DFFR_X1 my_filter_reg_samples_q_reg_12_ ( .D(my_filter_reg_samples_n32), 
        .CK(clk), .RN(my_filter_reg_samples_n46), .Q(my_filter_q_reg_samp_12_), 
        .QN(my_filter_reg_samples_n28) );
  DFFR_X1 my_filter_reg_samples_q_reg_13_ ( .D(my_filter_reg_samples_n31), 
        .CK(clk), .RN(my_filter_reg_samples_n46), .Q(my_filter_q_reg_samp_13_), 
        .QN(my_filter_reg_samples_n29) );
  CLKBUF_X1 my_filter_reg_coefficients_U352 ( .A(
        my_filter_reg_coefficients_n496), .Z(my_filter_reg_coefficients_n505)
         );
  CLKBUF_X1 my_filter_reg_coefficients_U351 ( .A(
        my_filter_reg_coefficients_n496), .Z(my_filter_reg_coefficients_n504)
         );
  CLKBUF_X1 my_filter_reg_coefficients_U350 ( .A(
        my_filter_reg_coefficients_n496), .Z(my_filter_reg_coefficients_n503)
         );
  CLKBUF_X1 my_filter_reg_coefficients_U349 ( .A(
        my_filter_reg_coefficients_n495), .Z(my_filter_reg_coefficients_n502)
         );
  CLKBUF_X1 my_filter_reg_coefficients_U348 ( .A(
        my_filter_reg_coefficients_n495), .Z(my_filter_reg_coefficients_n501)
         );
  CLKBUF_X1 my_filter_reg_coefficients_U347 ( .A(
        my_filter_reg_coefficients_n495), .Z(my_filter_reg_coefficients_n500)
         );
  CLKBUF_X1 my_filter_reg_coefficients_U346 ( .A(
        my_filter_reg_coefficients_n494), .Z(my_filter_reg_coefficients_n499)
         );
  CLKBUF_X1 my_filter_reg_coefficients_U345 ( .A(
        my_filter_reg_coefficients_n494), .Z(my_filter_reg_coefficients_n498)
         );
  CLKBUF_X1 my_filter_reg_coefficients_U344 ( .A(my_filter_n2), .Z(
        my_filter_reg_coefficients_n496) );
  CLKBUF_X1 my_filter_reg_coefficients_U343 ( .A(my_filter_n2), .Z(
        my_filter_reg_coefficients_n495) );
  CLKBUF_X1 my_filter_reg_coefficients_U342 ( .A(my_filter_n2), .Z(
        my_filter_reg_coefficients_n494) );
  INV_X1 my_filter_reg_coefficients_U341 ( .A(vin), .ZN(
        my_filter_reg_coefficients_n493) );
  NAND2_X1 my_filter_reg_coefficients_U340 ( .A1(
        my_filter_reg_coefficients_n482), .A2(b0[13]), .ZN(
        my_filter_reg_coefficients_n3) );
  OAI21_X1 my_filter_reg_coefficients_U339 ( .B1(
        my_filter_reg_coefficients_n480), .B2(my_filter_reg_coefficients_n286), 
        .A(my_filter_reg_coefficients_n3), .ZN(my_filter_reg_coefficients_n311) );
  NAND2_X1 my_filter_reg_coefficients_U338 ( .A1(b0[12]), .A2(
        my_filter_reg_coefficients_n492), .ZN(my_filter_reg_coefficients_n4)
         );
  OAI21_X1 my_filter_reg_coefficients_U337 ( .B1(
        my_filter_reg_coefficients_n480), .B2(my_filter_reg_coefficients_n285), 
        .A(my_filter_reg_coefficients_n4), .ZN(my_filter_reg_coefficients_n312) );
  NAND2_X1 my_filter_reg_coefficients_U336 ( .A1(b0[11]), .A2(
        my_filter_reg_coefficients_n491), .ZN(my_filter_reg_coefficients_n5)
         );
  OAI21_X1 my_filter_reg_coefficients_U335 ( .B1(
        my_filter_reg_coefficients_n480), .B2(my_filter_reg_coefficients_n284), 
        .A(my_filter_reg_coefficients_n5), .ZN(my_filter_reg_coefficients_n313) );
  NAND2_X1 my_filter_reg_coefficients_U334 ( .A1(b0[10]), .A2(
        my_filter_reg_coefficients_n490), .ZN(my_filter_reg_coefficients_n6)
         );
  OAI21_X1 my_filter_reg_coefficients_U333 ( .B1(
        my_filter_reg_coefficients_n480), .B2(my_filter_reg_coefficients_n283), 
        .A(my_filter_reg_coefficients_n6), .ZN(my_filter_reg_coefficients_n314) );
  NAND2_X1 my_filter_reg_coefficients_U332 ( .A1(b0[9]), .A2(
        my_filter_reg_coefficients_n489), .ZN(my_filter_reg_coefficients_n7)
         );
  OAI21_X1 my_filter_reg_coefficients_U331 ( .B1(
        my_filter_reg_coefficients_n480), .B2(my_filter_reg_coefficients_n282), 
        .A(my_filter_reg_coefficients_n7), .ZN(my_filter_reg_coefficients_n315) );
  NAND2_X1 my_filter_reg_coefficients_U330 ( .A1(b0[8]), .A2(
        my_filter_reg_coefficients_n488), .ZN(my_filter_reg_coefficients_n8)
         );
  OAI21_X1 my_filter_reg_coefficients_U329 ( .B1(
        my_filter_reg_coefficients_n480), .B2(my_filter_reg_coefficients_n281), 
        .A(my_filter_reg_coefficients_n8), .ZN(my_filter_reg_coefficients_n316) );
  NAND2_X1 my_filter_reg_coefficients_U328 ( .A1(b0[7]), .A2(
        my_filter_reg_coefficients_n487), .ZN(my_filter_reg_coefficients_n9)
         );
  OAI21_X1 my_filter_reg_coefficients_U327 ( .B1(
        my_filter_reg_coefficients_n480), .B2(my_filter_reg_coefficients_n280), 
        .A(my_filter_reg_coefficients_n9), .ZN(my_filter_reg_coefficients_n317) );
  NAND2_X1 my_filter_reg_coefficients_U326 ( .A1(b0[6]), .A2(
        my_filter_reg_coefficients_n486), .ZN(my_filter_reg_coefficients_n10)
         );
  OAI21_X1 my_filter_reg_coefficients_U325 ( .B1(
        my_filter_reg_coefficients_n480), .B2(my_filter_reg_coefficients_n279), 
        .A(my_filter_reg_coefficients_n10), .ZN(
        my_filter_reg_coefficients_n318) );
  NAND2_X1 my_filter_reg_coefficients_U324 ( .A1(b0[5]), .A2(
        my_filter_reg_coefficients_n485), .ZN(my_filter_reg_coefficients_n11)
         );
  OAI21_X1 my_filter_reg_coefficients_U323 ( .B1(
        my_filter_reg_coefficients_n480), .B2(my_filter_reg_coefficients_n278), 
        .A(my_filter_reg_coefficients_n11), .ZN(
        my_filter_reg_coefficients_n319) );
  NAND2_X1 my_filter_reg_coefficients_U322 ( .A1(b0[4]), .A2(
        my_filter_reg_coefficients_n481), .ZN(my_filter_reg_coefficients_n12)
         );
  OAI21_X1 my_filter_reg_coefficients_U321 ( .B1(
        my_filter_reg_coefficients_n480), .B2(my_filter_reg_coefficients_n277), 
        .A(my_filter_reg_coefficients_n12), .ZN(
        my_filter_reg_coefficients_n320) );
  NAND2_X1 my_filter_reg_coefficients_U320 ( .A1(b0[3]), .A2(
        my_filter_reg_coefficients_n492), .ZN(my_filter_reg_coefficients_n13)
         );
  OAI21_X1 my_filter_reg_coefficients_U319 ( .B1(
        my_filter_reg_coefficients_n479), .B2(my_filter_reg_coefficients_n276), 
        .A(my_filter_reg_coefficients_n13), .ZN(
        my_filter_reg_coefficients_n321) );
  NAND2_X1 my_filter_reg_coefficients_U318 ( .A1(b0[2]), .A2(
        my_filter_reg_coefficients_n492), .ZN(my_filter_reg_coefficients_n14)
         );
  OAI21_X1 my_filter_reg_coefficients_U317 ( .B1(
        my_filter_reg_coefficients_n479), .B2(my_filter_reg_coefficients_n275), 
        .A(my_filter_reg_coefficients_n14), .ZN(
        my_filter_reg_coefficients_n322) );
  NAND2_X1 my_filter_reg_coefficients_U316 ( .A1(b0[1]), .A2(
        my_filter_reg_coefficients_n492), .ZN(my_filter_reg_coefficients_n15)
         );
  OAI21_X1 my_filter_reg_coefficients_U315 ( .B1(
        my_filter_reg_coefficients_n479), .B2(my_filter_reg_coefficients_n274), 
        .A(my_filter_reg_coefficients_n15), .ZN(
        my_filter_reg_coefficients_n323) );
  NAND2_X1 my_filter_reg_coefficients_U314 ( .A1(b0[0]), .A2(
        my_filter_reg_coefficients_n492), .ZN(my_filter_reg_coefficients_n16)
         );
  OAI21_X1 my_filter_reg_coefficients_U313 ( .B1(
        my_filter_reg_coefficients_n479), .B2(my_filter_reg_coefficients_n273), 
        .A(my_filter_reg_coefficients_n16), .ZN(
        my_filter_reg_coefficients_n324) );
  NAND2_X1 my_filter_reg_coefficients_U312 ( .A1(b1[13]), .A2(
        my_filter_reg_coefficients_n492), .ZN(my_filter_reg_coefficients_n17)
         );
  OAI21_X1 my_filter_reg_coefficients_U311 ( .B1(
        my_filter_reg_coefficients_n479), .B2(my_filter_reg_coefficients_n272), 
        .A(my_filter_reg_coefficients_n17), .ZN(
        my_filter_reg_coefficients_n325) );
  NAND2_X1 my_filter_reg_coefficients_U310 ( .A1(b1[12]), .A2(
        my_filter_reg_coefficients_n492), .ZN(my_filter_reg_coefficients_n18)
         );
  OAI21_X1 my_filter_reg_coefficients_U309 ( .B1(
        my_filter_reg_coefficients_n479), .B2(my_filter_reg_coefficients_n271), 
        .A(my_filter_reg_coefficients_n18), .ZN(
        my_filter_reg_coefficients_n326) );
  NAND2_X1 my_filter_reg_coefficients_U308 ( .A1(b1[11]), .A2(
        my_filter_reg_coefficients_n492), .ZN(my_filter_reg_coefficients_n19)
         );
  OAI21_X1 my_filter_reg_coefficients_U307 ( .B1(
        my_filter_reg_coefficients_n479), .B2(my_filter_reg_coefficients_n270), 
        .A(my_filter_reg_coefficients_n19), .ZN(
        my_filter_reg_coefficients_n327) );
  NAND2_X1 my_filter_reg_coefficients_U306 ( .A1(b1[10]), .A2(
        my_filter_reg_coefficients_n492), .ZN(my_filter_reg_coefficients_n20)
         );
  OAI21_X1 my_filter_reg_coefficients_U305 ( .B1(
        my_filter_reg_coefficients_n479), .B2(my_filter_reg_coefficients_n269), 
        .A(my_filter_reg_coefficients_n20), .ZN(
        my_filter_reg_coefficients_n328) );
  NAND2_X1 my_filter_reg_coefficients_U304 ( .A1(b1[9]), .A2(
        my_filter_reg_coefficients_n492), .ZN(my_filter_reg_coefficients_n21)
         );
  OAI21_X1 my_filter_reg_coefficients_U303 ( .B1(
        my_filter_reg_coefficients_n479), .B2(my_filter_reg_coefficients_n268), 
        .A(my_filter_reg_coefficients_n21), .ZN(
        my_filter_reg_coefficients_n329) );
  NAND2_X1 my_filter_reg_coefficients_U302 ( .A1(b1[8]), .A2(
        my_filter_reg_coefficients_n492), .ZN(my_filter_reg_coefficients_n22)
         );
  OAI21_X1 my_filter_reg_coefficients_U301 ( .B1(
        my_filter_reg_coefficients_n479), .B2(my_filter_reg_coefficients_n267), 
        .A(my_filter_reg_coefficients_n22), .ZN(
        my_filter_reg_coefficients_n330) );
  NAND2_X1 my_filter_reg_coefficients_U300 ( .A1(b1[7]), .A2(
        my_filter_reg_coefficients_n492), .ZN(my_filter_reg_coefficients_n23)
         );
  OAI21_X1 my_filter_reg_coefficients_U299 ( .B1(
        my_filter_reg_coefficients_n479), .B2(my_filter_reg_coefficients_n266), 
        .A(my_filter_reg_coefficients_n23), .ZN(
        my_filter_reg_coefficients_n331) );
  NAND2_X1 my_filter_reg_coefficients_U298 ( .A1(b1[6]), .A2(
        my_filter_reg_coefficients_n492), .ZN(my_filter_reg_coefficients_n24)
         );
  OAI21_X1 my_filter_reg_coefficients_U297 ( .B1(
        my_filter_reg_coefficients_n479), .B2(my_filter_reg_coefficients_n265), 
        .A(my_filter_reg_coefficients_n24), .ZN(
        my_filter_reg_coefficients_n332) );
  NAND2_X1 my_filter_reg_coefficients_U296 ( .A1(b1[5]), .A2(
        my_filter_reg_coefficients_n491), .ZN(my_filter_reg_coefficients_n25)
         );
  OAI21_X1 my_filter_reg_coefficients_U295 ( .B1(
        my_filter_reg_coefficients_n478), .B2(my_filter_reg_coefficients_n264), 
        .A(my_filter_reg_coefficients_n25), .ZN(
        my_filter_reg_coefficients_n333) );
  NAND2_X1 my_filter_reg_coefficients_U294 ( .A1(b1[4]), .A2(
        my_filter_reg_coefficients_n491), .ZN(my_filter_reg_coefficients_n26)
         );
  OAI21_X1 my_filter_reg_coefficients_U293 ( .B1(
        my_filter_reg_coefficients_n478), .B2(my_filter_reg_coefficients_n263), 
        .A(my_filter_reg_coefficients_n26), .ZN(
        my_filter_reg_coefficients_n334) );
  NAND2_X1 my_filter_reg_coefficients_U292 ( .A1(b1[3]), .A2(
        my_filter_reg_coefficients_n491), .ZN(my_filter_reg_coefficients_n27)
         );
  OAI21_X1 my_filter_reg_coefficients_U291 ( .B1(
        my_filter_reg_coefficients_n478), .B2(my_filter_reg_coefficients_n262), 
        .A(my_filter_reg_coefficients_n27), .ZN(
        my_filter_reg_coefficients_n335) );
  NAND2_X1 my_filter_reg_coefficients_U290 ( .A1(b1[2]), .A2(
        my_filter_reg_coefficients_n491), .ZN(my_filter_reg_coefficients_n28)
         );
  OAI21_X1 my_filter_reg_coefficients_U289 ( .B1(
        my_filter_reg_coefficients_n478), .B2(my_filter_reg_coefficients_n261), 
        .A(my_filter_reg_coefficients_n28), .ZN(
        my_filter_reg_coefficients_n336) );
  NAND2_X1 my_filter_reg_coefficients_U288 ( .A1(b1[1]), .A2(
        my_filter_reg_coefficients_n491), .ZN(my_filter_reg_coefficients_n29)
         );
  OAI21_X1 my_filter_reg_coefficients_U287 ( .B1(
        my_filter_reg_coefficients_n478), .B2(my_filter_reg_coefficients_n260), 
        .A(my_filter_reg_coefficients_n29), .ZN(
        my_filter_reg_coefficients_n337) );
  NAND2_X1 my_filter_reg_coefficients_U286 ( .A1(b1[0]), .A2(
        my_filter_reg_coefficients_n491), .ZN(my_filter_reg_coefficients_n30)
         );
  OAI21_X1 my_filter_reg_coefficients_U285 ( .B1(
        my_filter_reg_coefficients_n478), .B2(my_filter_reg_coefficients_n259), 
        .A(my_filter_reg_coefficients_n30), .ZN(
        my_filter_reg_coefficients_n338) );
  NAND2_X1 my_filter_reg_coefficients_U284 ( .A1(b2[13]), .A2(
        my_filter_reg_coefficients_n491), .ZN(my_filter_reg_coefficients_n31)
         );
  OAI21_X1 my_filter_reg_coefficients_U283 ( .B1(
        my_filter_reg_coefficients_n478), .B2(my_filter_reg_coefficients_n258), 
        .A(my_filter_reg_coefficients_n31), .ZN(
        my_filter_reg_coefficients_n339) );
  NAND2_X1 my_filter_reg_coefficients_U282 ( .A1(b2[12]), .A2(
        my_filter_reg_coefficients_n491), .ZN(my_filter_reg_coefficients_n32)
         );
  OAI21_X1 my_filter_reg_coefficients_U281 ( .B1(
        my_filter_reg_coefficients_n478), .B2(my_filter_reg_coefficients_n257), 
        .A(my_filter_reg_coefficients_n32), .ZN(
        my_filter_reg_coefficients_n340) );
  NAND2_X1 my_filter_reg_coefficients_U280 ( .A1(b2[11]), .A2(
        my_filter_reg_coefficients_n491), .ZN(my_filter_reg_coefficients_n33)
         );
  OAI21_X1 my_filter_reg_coefficients_U279 ( .B1(
        my_filter_reg_coefficients_n478), .B2(my_filter_reg_coefficients_n256), 
        .A(my_filter_reg_coefficients_n33), .ZN(
        my_filter_reg_coefficients_n341) );
  NAND2_X1 my_filter_reg_coefficients_U278 ( .A1(b2[10]), .A2(
        my_filter_reg_coefficients_n491), .ZN(my_filter_reg_coefficients_n34)
         );
  OAI21_X1 my_filter_reg_coefficients_U277 ( .B1(
        my_filter_reg_coefficients_n478), .B2(my_filter_reg_coefficients_n255), 
        .A(my_filter_reg_coefficients_n34), .ZN(
        my_filter_reg_coefficients_n342) );
  NAND2_X1 my_filter_reg_coefficients_U276 ( .A1(b2[9]), .A2(
        my_filter_reg_coefficients_n491), .ZN(my_filter_reg_coefficients_n35)
         );
  OAI21_X1 my_filter_reg_coefficients_U275 ( .B1(
        my_filter_reg_coefficients_n478), .B2(my_filter_reg_coefficients_n254), 
        .A(my_filter_reg_coefficients_n35), .ZN(
        my_filter_reg_coefficients_n343) );
  NAND2_X1 my_filter_reg_coefficients_U274 ( .A1(b2[8]), .A2(
        my_filter_reg_coefficients_n491), .ZN(my_filter_reg_coefficients_n36)
         );
  OAI21_X1 my_filter_reg_coefficients_U273 ( .B1(
        my_filter_reg_coefficients_n478), .B2(my_filter_reg_coefficients_n253), 
        .A(my_filter_reg_coefficients_n36), .ZN(
        my_filter_reg_coefficients_n344) );
  NAND2_X1 my_filter_reg_coefficients_U272 ( .A1(b2[7]), .A2(
        my_filter_reg_coefficients_n490), .ZN(my_filter_reg_coefficients_n37)
         );
  OAI21_X1 my_filter_reg_coefficients_U271 ( .B1(
        my_filter_reg_coefficients_n477), .B2(my_filter_reg_coefficients_n252), 
        .A(my_filter_reg_coefficients_n37), .ZN(
        my_filter_reg_coefficients_n345) );
  NAND2_X1 my_filter_reg_coefficients_U270 ( .A1(b2[6]), .A2(
        my_filter_reg_coefficients_n490), .ZN(my_filter_reg_coefficients_n38)
         );
  OAI21_X1 my_filter_reg_coefficients_U269 ( .B1(
        my_filter_reg_coefficients_n477), .B2(my_filter_reg_coefficients_n251), 
        .A(my_filter_reg_coefficients_n38), .ZN(
        my_filter_reg_coefficients_n346) );
  NAND2_X1 my_filter_reg_coefficients_U268 ( .A1(b2[5]), .A2(
        my_filter_reg_coefficients_n490), .ZN(my_filter_reg_coefficients_n39)
         );
  OAI21_X1 my_filter_reg_coefficients_U267 ( .B1(
        my_filter_reg_coefficients_n477), .B2(my_filter_reg_coefficients_n250), 
        .A(my_filter_reg_coefficients_n39), .ZN(
        my_filter_reg_coefficients_n347) );
  NAND2_X1 my_filter_reg_coefficients_U266 ( .A1(b2[4]), .A2(
        my_filter_reg_coefficients_n490), .ZN(my_filter_reg_coefficients_n40)
         );
  OAI21_X1 my_filter_reg_coefficients_U265 ( .B1(
        my_filter_reg_coefficients_n477), .B2(my_filter_reg_coefficients_n249), 
        .A(my_filter_reg_coefficients_n40), .ZN(
        my_filter_reg_coefficients_n348) );
  NAND2_X1 my_filter_reg_coefficients_U264 ( .A1(b2[3]), .A2(
        my_filter_reg_coefficients_n490), .ZN(my_filter_reg_coefficients_n41)
         );
  OAI21_X1 my_filter_reg_coefficients_U263 ( .B1(
        my_filter_reg_coefficients_n477), .B2(my_filter_reg_coefficients_n248), 
        .A(my_filter_reg_coefficients_n41), .ZN(
        my_filter_reg_coefficients_n349) );
  NAND2_X1 my_filter_reg_coefficients_U262 ( .A1(b2[2]), .A2(
        my_filter_reg_coefficients_n490), .ZN(my_filter_reg_coefficients_n42)
         );
  OAI21_X1 my_filter_reg_coefficients_U261 ( .B1(
        my_filter_reg_coefficients_n477), .B2(my_filter_reg_coefficients_n247), 
        .A(my_filter_reg_coefficients_n42), .ZN(
        my_filter_reg_coefficients_n350) );
  NAND2_X1 my_filter_reg_coefficients_U260 ( .A1(b2[1]), .A2(
        my_filter_reg_coefficients_n490), .ZN(my_filter_reg_coefficients_n43)
         );
  OAI21_X1 my_filter_reg_coefficients_U259 ( .B1(
        my_filter_reg_coefficients_n477), .B2(my_filter_reg_coefficients_n246), 
        .A(my_filter_reg_coefficients_n43), .ZN(
        my_filter_reg_coefficients_n351) );
  NAND2_X1 my_filter_reg_coefficients_U258 ( .A1(b2[0]), .A2(
        my_filter_reg_coefficients_n490), .ZN(my_filter_reg_coefficients_n44)
         );
  OAI21_X1 my_filter_reg_coefficients_U257 ( .B1(
        my_filter_reg_coefficients_n477), .B2(my_filter_reg_coefficients_n245), 
        .A(my_filter_reg_coefficients_n44), .ZN(
        my_filter_reg_coefficients_n352) );
  NAND2_X1 my_filter_reg_coefficients_U256 ( .A1(b3[13]), .A2(
        my_filter_reg_coefficients_n490), .ZN(my_filter_reg_coefficients_n45)
         );
  OAI21_X1 my_filter_reg_coefficients_U255 ( .B1(
        my_filter_reg_coefficients_n477), .B2(my_filter_reg_coefficients_n244), 
        .A(my_filter_reg_coefficients_n45), .ZN(
        my_filter_reg_coefficients_n353) );
  NAND2_X1 my_filter_reg_coefficients_U254 ( .A1(b3[12]), .A2(
        my_filter_reg_coefficients_n490), .ZN(my_filter_reg_coefficients_n46)
         );
  OAI21_X1 my_filter_reg_coefficients_U253 ( .B1(
        my_filter_reg_coefficients_n477), .B2(my_filter_reg_coefficients_n243), 
        .A(my_filter_reg_coefficients_n46), .ZN(
        my_filter_reg_coefficients_n354) );
  NAND2_X1 my_filter_reg_coefficients_U252 ( .A1(b3[11]), .A2(
        my_filter_reg_coefficients_n490), .ZN(my_filter_reg_coefficients_n47)
         );
  OAI21_X1 my_filter_reg_coefficients_U251 ( .B1(
        my_filter_reg_coefficients_n477), .B2(my_filter_reg_coefficients_n242), 
        .A(my_filter_reg_coefficients_n47), .ZN(
        my_filter_reg_coefficients_n355) );
  NAND2_X1 my_filter_reg_coefficients_U250 ( .A1(b3[10]), .A2(
        my_filter_reg_coefficients_n490), .ZN(my_filter_reg_coefficients_n48)
         );
  OAI21_X1 my_filter_reg_coefficients_U249 ( .B1(
        my_filter_reg_coefficients_n477), .B2(my_filter_reg_coefficients_n241), 
        .A(my_filter_reg_coefficients_n48), .ZN(
        my_filter_reg_coefficients_n356) );
  NAND2_X1 my_filter_reg_coefficients_U248 ( .A1(b3[9]), .A2(
        my_filter_reg_coefficients_n489), .ZN(my_filter_reg_coefficients_n49)
         );
  OAI21_X1 my_filter_reg_coefficients_U247 ( .B1(
        my_filter_reg_coefficients_n476), .B2(my_filter_reg_coefficients_n240), 
        .A(my_filter_reg_coefficients_n49), .ZN(
        my_filter_reg_coefficients_n357) );
  NAND2_X1 my_filter_reg_coefficients_U246 ( .A1(b3[8]), .A2(
        my_filter_reg_coefficients_n489), .ZN(my_filter_reg_coefficients_n50)
         );
  OAI21_X1 my_filter_reg_coefficients_U245 ( .B1(
        my_filter_reg_coefficients_n476), .B2(my_filter_reg_coefficients_n239), 
        .A(my_filter_reg_coefficients_n50), .ZN(
        my_filter_reg_coefficients_n358) );
  NAND2_X1 my_filter_reg_coefficients_U244 ( .A1(b3[7]), .A2(
        my_filter_reg_coefficients_n489), .ZN(my_filter_reg_coefficients_n51)
         );
  OAI21_X1 my_filter_reg_coefficients_U243 ( .B1(
        my_filter_reg_coefficients_n476), .B2(my_filter_reg_coefficients_n238), 
        .A(my_filter_reg_coefficients_n51), .ZN(
        my_filter_reg_coefficients_n359) );
  NAND2_X1 my_filter_reg_coefficients_U242 ( .A1(b3[6]), .A2(
        my_filter_reg_coefficients_n489), .ZN(my_filter_reg_coefficients_n52)
         );
  OAI21_X1 my_filter_reg_coefficients_U241 ( .B1(
        my_filter_reg_coefficients_n476), .B2(my_filter_reg_coefficients_n237), 
        .A(my_filter_reg_coefficients_n52), .ZN(
        my_filter_reg_coefficients_n360) );
  NAND2_X1 my_filter_reg_coefficients_U240 ( .A1(b3[5]), .A2(
        my_filter_reg_coefficients_n489), .ZN(my_filter_reg_coefficients_n53)
         );
  OAI21_X1 my_filter_reg_coefficients_U239 ( .B1(
        my_filter_reg_coefficients_n476), .B2(my_filter_reg_coefficients_n236), 
        .A(my_filter_reg_coefficients_n53), .ZN(
        my_filter_reg_coefficients_n361) );
  NAND2_X1 my_filter_reg_coefficients_U238 ( .A1(b3[4]), .A2(
        my_filter_reg_coefficients_n489), .ZN(my_filter_reg_coefficients_n54)
         );
  OAI21_X1 my_filter_reg_coefficients_U237 ( .B1(
        my_filter_reg_coefficients_n476), .B2(my_filter_reg_coefficients_n235), 
        .A(my_filter_reg_coefficients_n54), .ZN(
        my_filter_reg_coefficients_n362) );
  NAND2_X1 my_filter_reg_coefficients_U236 ( .A1(b3[3]), .A2(
        my_filter_reg_coefficients_n489), .ZN(my_filter_reg_coefficients_n55)
         );
  OAI21_X1 my_filter_reg_coefficients_U235 ( .B1(
        my_filter_reg_coefficients_n476), .B2(my_filter_reg_coefficients_n234), 
        .A(my_filter_reg_coefficients_n55), .ZN(
        my_filter_reg_coefficients_n363) );
  NAND2_X1 my_filter_reg_coefficients_U234 ( .A1(b3[2]), .A2(
        my_filter_reg_coefficients_n489), .ZN(my_filter_reg_coefficients_n56)
         );
  OAI21_X1 my_filter_reg_coefficients_U233 ( .B1(
        my_filter_reg_coefficients_n476), .B2(my_filter_reg_coefficients_n233), 
        .A(my_filter_reg_coefficients_n56), .ZN(
        my_filter_reg_coefficients_n364) );
  NAND2_X1 my_filter_reg_coefficients_U232 ( .A1(b3[1]), .A2(
        my_filter_reg_coefficients_n489), .ZN(my_filter_reg_coefficients_n57)
         );
  OAI21_X1 my_filter_reg_coefficients_U231 ( .B1(
        my_filter_reg_coefficients_n476), .B2(my_filter_reg_coefficients_n232), 
        .A(my_filter_reg_coefficients_n57), .ZN(
        my_filter_reg_coefficients_n365) );
  NAND2_X1 my_filter_reg_coefficients_U230 ( .A1(b3[0]), .A2(
        my_filter_reg_coefficients_n489), .ZN(my_filter_reg_coefficients_n58)
         );
  OAI21_X1 my_filter_reg_coefficients_U229 ( .B1(
        my_filter_reg_coefficients_n476), .B2(my_filter_reg_coefficients_n231), 
        .A(my_filter_reg_coefficients_n58), .ZN(
        my_filter_reg_coefficients_n366) );
  NAND2_X1 my_filter_reg_coefficients_U228 ( .A1(b4[13]), .A2(
        my_filter_reg_coefficients_n489), .ZN(my_filter_reg_coefficients_n59)
         );
  OAI21_X1 my_filter_reg_coefficients_U227 ( .B1(
        my_filter_reg_coefficients_n476), .B2(my_filter_reg_coefficients_n230), 
        .A(my_filter_reg_coefficients_n59), .ZN(
        my_filter_reg_coefficients_n367) );
  NAND2_X1 my_filter_reg_coefficients_U226 ( .A1(b4[12]), .A2(
        my_filter_reg_coefficients_n489), .ZN(my_filter_reg_coefficients_n60)
         );
  OAI21_X1 my_filter_reg_coefficients_U225 ( .B1(
        my_filter_reg_coefficients_n476), .B2(my_filter_reg_coefficients_n229), 
        .A(my_filter_reg_coefficients_n60), .ZN(
        my_filter_reg_coefficients_n368) );
  NAND2_X1 my_filter_reg_coefficients_U224 ( .A1(b4[11]), .A2(
        my_filter_reg_coefficients_n488), .ZN(my_filter_reg_coefficients_n61)
         );
  OAI21_X1 my_filter_reg_coefficients_U223 ( .B1(
        my_filter_reg_coefficients_n475), .B2(my_filter_reg_coefficients_n228), 
        .A(my_filter_reg_coefficients_n61), .ZN(
        my_filter_reg_coefficients_n369) );
  NAND2_X1 my_filter_reg_coefficients_U222 ( .A1(b4[10]), .A2(
        my_filter_reg_coefficients_n488), .ZN(my_filter_reg_coefficients_n62)
         );
  OAI21_X1 my_filter_reg_coefficients_U221 ( .B1(
        my_filter_reg_coefficients_n475), .B2(my_filter_reg_coefficients_n227), 
        .A(my_filter_reg_coefficients_n62), .ZN(
        my_filter_reg_coefficients_n370) );
  NAND2_X1 my_filter_reg_coefficients_U220 ( .A1(b4[9]), .A2(
        my_filter_reg_coefficients_n488), .ZN(my_filter_reg_coefficients_n63)
         );
  OAI21_X1 my_filter_reg_coefficients_U219 ( .B1(
        my_filter_reg_coefficients_n475), .B2(my_filter_reg_coefficients_n226), 
        .A(my_filter_reg_coefficients_n63), .ZN(
        my_filter_reg_coefficients_n371) );
  NAND2_X1 my_filter_reg_coefficients_U218 ( .A1(b4[8]), .A2(
        my_filter_reg_coefficients_n488), .ZN(my_filter_reg_coefficients_n64)
         );
  OAI21_X1 my_filter_reg_coefficients_U217 ( .B1(
        my_filter_reg_coefficients_n475), .B2(my_filter_reg_coefficients_n225), 
        .A(my_filter_reg_coefficients_n64), .ZN(
        my_filter_reg_coefficients_n372) );
  NAND2_X1 my_filter_reg_coefficients_U216 ( .A1(b4[7]), .A2(
        my_filter_reg_coefficients_n488), .ZN(my_filter_reg_coefficients_n65)
         );
  OAI21_X1 my_filter_reg_coefficients_U215 ( .B1(
        my_filter_reg_coefficients_n475), .B2(my_filter_reg_coefficients_n224), 
        .A(my_filter_reg_coefficients_n65), .ZN(
        my_filter_reg_coefficients_n373) );
  NAND2_X1 my_filter_reg_coefficients_U214 ( .A1(b4[6]), .A2(
        my_filter_reg_coefficients_n488), .ZN(my_filter_reg_coefficients_n66)
         );
  OAI21_X1 my_filter_reg_coefficients_U213 ( .B1(
        my_filter_reg_coefficients_n475), .B2(my_filter_reg_coefficients_n223), 
        .A(my_filter_reg_coefficients_n66), .ZN(
        my_filter_reg_coefficients_n374) );
  NAND2_X1 my_filter_reg_coefficients_U212 ( .A1(b4[5]), .A2(
        my_filter_reg_coefficients_n488), .ZN(my_filter_reg_coefficients_n67)
         );
  OAI21_X1 my_filter_reg_coefficients_U211 ( .B1(
        my_filter_reg_coefficients_n475), .B2(my_filter_reg_coefficients_n222), 
        .A(my_filter_reg_coefficients_n67), .ZN(
        my_filter_reg_coefficients_n375) );
  NAND2_X1 my_filter_reg_coefficients_U210 ( .A1(b4[4]), .A2(
        my_filter_reg_coefficients_n488), .ZN(my_filter_reg_coefficients_n68)
         );
  OAI21_X1 my_filter_reg_coefficients_U209 ( .B1(
        my_filter_reg_coefficients_n475), .B2(my_filter_reg_coefficients_n221), 
        .A(my_filter_reg_coefficients_n68), .ZN(
        my_filter_reg_coefficients_n376) );
  NAND2_X1 my_filter_reg_coefficients_U208 ( .A1(b4[3]), .A2(
        my_filter_reg_coefficients_n488), .ZN(my_filter_reg_coefficients_n69)
         );
  OAI21_X1 my_filter_reg_coefficients_U207 ( .B1(
        my_filter_reg_coefficients_n475), .B2(my_filter_reg_coefficients_n220), 
        .A(my_filter_reg_coefficients_n69), .ZN(
        my_filter_reg_coefficients_n377) );
  NAND2_X1 my_filter_reg_coefficients_U206 ( .A1(b4[2]), .A2(
        my_filter_reg_coefficients_n488), .ZN(my_filter_reg_coefficients_n70)
         );
  OAI21_X1 my_filter_reg_coefficients_U205 ( .B1(
        my_filter_reg_coefficients_n475), .B2(my_filter_reg_coefficients_n219), 
        .A(my_filter_reg_coefficients_n70), .ZN(
        my_filter_reg_coefficients_n378) );
  NAND2_X1 my_filter_reg_coefficients_U204 ( .A1(b4[1]), .A2(
        my_filter_reg_coefficients_n488), .ZN(my_filter_reg_coefficients_n71)
         );
  OAI21_X1 my_filter_reg_coefficients_U203 ( .B1(
        my_filter_reg_coefficients_n475), .B2(my_filter_reg_coefficients_n218), 
        .A(my_filter_reg_coefficients_n71), .ZN(
        my_filter_reg_coefficients_n379) );
  NAND2_X1 my_filter_reg_coefficients_U202 ( .A1(b4[0]), .A2(
        my_filter_reg_coefficients_n488), .ZN(my_filter_reg_coefficients_n72)
         );
  OAI21_X1 my_filter_reg_coefficients_U201 ( .B1(
        my_filter_reg_coefficients_n475), .B2(my_filter_reg_coefficients_n217), 
        .A(my_filter_reg_coefficients_n72), .ZN(
        my_filter_reg_coefficients_n380) );
  NAND2_X1 my_filter_reg_coefficients_U200 ( .A1(b5[13]), .A2(
        my_filter_reg_coefficients_n487), .ZN(my_filter_reg_coefficients_n73)
         );
  OAI21_X1 my_filter_reg_coefficients_U199 ( .B1(
        my_filter_reg_coefficients_n474), .B2(my_filter_reg_coefficients_n216), 
        .A(my_filter_reg_coefficients_n73), .ZN(
        my_filter_reg_coefficients_n381) );
  NAND2_X1 my_filter_reg_coefficients_U198 ( .A1(b5[12]), .A2(
        my_filter_reg_coefficients_n487), .ZN(my_filter_reg_coefficients_n74)
         );
  OAI21_X1 my_filter_reg_coefficients_U197 ( .B1(
        my_filter_reg_coefficients_n474), .B2(my_filter_reg_coefficients_n215), 
        .A(my_filter_reg_coefficients_n74), .ZN(
        my_filter_reg_coefficients_n382) );
  NAND2_X1 my_filter_reg_coefficients_U196 ( .A1(b5[11]), .A2(
        my_filter_reg_coefficients_n487), .ZN(my_filter_reg_coefficients_n75)
         );
  OAI21_X1 my_filter_reg_coefficients_U195 ( .B1(
        my_filter_reg_coefficients_n474), .B2(my_filter_reg_coefficients_n214), 
        .A(my_filter_reg_coefficients_n75), .ZN(
        my_filter_reg_coefficients_n383) );
  NAND2_X1 my_filter_reg_coefficients_U194 ( .A1(b5[10]), .A2(
        my_filter_reg_coefficients_n487), .ZN(my_filter_reg_coefficients_n76)
         );
  OAI21_X1 my_filter_reg_coefficients_U193 ( .B1(
        my_filter_reg_coefficients_n474), .B2(my_filter_reg_coefficients_n213), 
        .A(my_filter_reg_coefficients_n76), .ZN(
        my_filter_reg_coefficients_n384) );
  NAND2_X1 my_filter_reg_coefficients_U192 ( .A1(b5[9]), .A2(
        my_filter_reg_coefficients_n487), .ZN(my_filter_reg_coefficients_n77)
         );
  OAI21_X1 my_filter_reg_coefficients_U191 ( .B1(
        my_filter_reg_coefficients_n474), .B2(my_filter_reg_coefficients_n212), 
        .A(my_filter_reg_coefficients_n77), .ZN(
        my_filter_reg_coefficients_n385) );
  NAND2_X1 my_filter_reg_coefficients_U190 ( .A1(b5[8]), .A2(
        my_filter_reg_coefficients_n487), .ZN(my_filter_reg_coefficients_n78)
         );
  OAI21_X1 my_filter_reg_coefficients_U189 ( .B1(
        my_filter_reg_coefficients_n474), .B2(my_filter_reg_coefficients_n211), 
        .A(my_filter_reg_coefficients_n78), .ZN(
        my_filter_reg_coefficients_n386) );
  NAND2_X1 my_filter_reg_coefficients_U188 ( .A1(b5[7]), .A2(
        my_filter_reg_coefficients_n487), .ZN(my_filter_reg_coefficients_n79)
         );
  OAI21_X1 my_filter_reg_coefficients_U187 ( .B1(
        my_filter_reg_coefficients_n474), .B2(my_filter_reg_coefficients_n210), 
        .A(my_filter_reg_coefficients_n79), .ZN(
        my_filter_reg_coefficients_n387) );
  NAND2_X1 my_filter_reg_coefficients_U186 ( .A1(b5[6]), .A2(
        my_filter_reg_coefficients_n487), .ZN(my_filter_reg_coefficients_n80)
         );
  OAI21_X1 my_filter_reg_coefficients_U185 ( .B1(
        my_filter_reg_coefficients_n474), .B2(my_filter_reg_coefficients_n209), 
        .A(my_filter_reg_coefficients_n80), .ZN(
        my_filter_reg_coefficients_n388) );
  NAND2_X1 my_filter_reg_coefficients_U184 ( .A1(b5[5]), .A2(
        my_filter_reg_coefficients_n487), .ZN(my_filter_reg_coefficients_n81)
         );
  OAI21_X1 my_filter_reg_coefficients_U183 ( .B1(
        my_filter_reg_coefficients_n474), .B2(my_filter_reg_coefficients_n208), 
        .A(my_filter_reg_coefficients_n81), .ZN(
        my_filter_reg_coefficients_n389) );
  NAND2_X1 my_filter_reg_coefficients_U182 ( .A1(b5[4]), .A2(
        my_filter_reg_coefficients_n487), .ZN(my_filter_reg_coefficients_n82)
         );
  OAI21_X1 my_filter_reg_coefficients_U181 ( .B1(
        my_filter_reg_coefficients_n474), .B2(my_filter_reg_coefficients_n207), 
        .A(my_filter_reg_coefficients_n82), .ZN(
        my_filter_reg_coefficients_n390) );
  NAND2_X1 my_filter_reg_coefficients_U180 ( .A1(b5[3]), .A2(
        my_filter_reg_coefficients_n487), .ZN(my_filter_reg_coefficients_n83)
         );
  OAI21_X1 my_filter_reg_coefficients_U179 ( .B1(
        my_filter_reg_coefficients_n474), .B2(my_filter_reg_coefficients_n206), 
        .A(my_filter_reg_coefficients_n83), .ZN(
        my_filter_reg_coefficients_n391) );
  NAND2_X1 my_filter_reg_coefficients_U178 ( .A1(b5[2]), .A2(
        my_filter_reg_coefficients_n487), .ZN(my_filter_reg_coefficients_n84)
         );
  OAI21_X1 my_filter_reg_coefficients_U177 ( .B1(
        my_filter_reg_coefficients_n474), .B2(my_filter_reg_coefficients_n205), 
        .A(my_filter_reg_coefficients_n84), .ZN(
        my_filter_reg_coefficients_n392) );
  NAND2_X1 my_filter_reg_coefficients_U176 ( .A1(b5[1]), .A2(
        my_filter_reg_coefficients_n486), .ZN(my_filter_reg_coefficients_n85)
         );
  OAI21_X1 my_filter_reg_coefficients_U175 ( .B1(
        my_filter_reg_coefficients_n473), .B2(my_filter_reg_coefficients_n204), 
        .A(my_filter_reg_coefficients_n85), .ZN(
        my_filter_reg_coefficients_n393) );
  NAND2_X1 my_filter_reg_coefficients_U174 ( .A1(b5[0]), .A2(
        my_filter_reg_coefficients_n486), .ZN(my_filter_reg_coefficients_n86)
         );
  OAI21_X1 my_filter_reg_coefficients_U173 ( .B1(
        my_filter_reg_coefficients_n473), .B2(my_filter_reg_coefficients_n203), 
        .A(my_filter_reg_coefficients_n86), .ZN(
        my_filter_reg_coefficients_n394) );
  NAND2_X1 my_filter_reg_coefficients_U172 ( .A1(b6[13]), .A2(
        my_filter_reg_coefficients_n486), .ZN(my_filter_reg_coefficients_n87)
         );
  OAI21_X1 my_filter_reg_coefficients_U171 ( .B1(
        my_filter_reg_coefficients_n473), .B2(my_filter_reg_coefficients_n202), 
        .A(my_filter_reg_coefficients_n87), .ZN(
        my_filter_reg_coefficients_n395) );
  NAND2_X1 my_filter_reg_coefficients_U170 ( .A1(b6[12]), .A2(
        my_filter_reg_coefficients_n486), .ZN(my_filter_reg_coefficients_n88)
         );
  OAI21_X1 my_filter_reg_coefficients_U169 ( .B1(
        my_filter_reg_coefficients_n473), .B2(my_filter_reg_coefficients_n201), 
        .A(my_filter_reg_coefficients_n88), .ZN(
        my_filter_reg_coefficients_n396) );
  NAND2_X1 my_filter_reg_coefficients_U168 ( .A1(b6[11]), .A2(
        my_filter_reg_coefficients_n486), .ZN(my_filter_reg_coefficients_n89)
         );
  OAI21_X1 my_filter_reg_coefficients_U167 ( .B1(
        my_filter_reg_coefficients_n473), .B2(my_filter_reg_coefficients_n200), 
        .A(my_filter_reg_coefficients_n89), .ZN(
        my_filter_reg_coefficients_n397) );
  NAND2_X1 my_filter_reg_coefficients_U166 ( .A1(b6[10]), .A2(
        my_filter_reg_coefficients_n486), .ZN(my_filter_reg_coefficients_n90)
         );
  OAI21_X1 my_filter_reg_coefficients_U165 ( .B1(
        my_filter_reg_coefficients_n473), .B2(my_filter_reg_coefficients_n199), 
        .A(my_filter_reg_coefficients_n90), .ZN(
        my_filter_reg_coefficients_n398) );
  NAND2_X1 my_filter_reg_coefficients_U164 ( .A1(b6[9]), .A2(
        my_filter_reg_coefficients_n486), .ZN(my_filter_reg_coefficients_n91)
         );
  OAI21_X1 my_filter_reg_coefficients_U163 ( .B1(
        my_filter_reg_coefficients_n473), .B2(my_filter_reg_coefficients_n198), 
        .A(my_filter_reg_coefficients_n91), .ZN(
        my_filter_reg_coefficients_n399) );
  NAND2_X1 my_filter_reg_coefficients_U162 ( .A1(b6[8]), .A2(
        my_filter_reg_coefficients_n486), .ZN(my_filter_reg_coefficients_n92)
         );
  OAI21_X1 my_filter_reg_coefficients_U161 ( .B1(
        my_filter_reg_coefficients_n473), .B2(my_filter_reg_coefficients_n197), 
        .A(my_filter_reg_coefficients_n92), .ZN(
        my_filter_reg_coefficients_n400) );
  NAND2_X1 my_filter_reg_coefficients_U160 ( .A1(b6[7]), .A2(
        my_filter_reg_coefficients_n486), .ZN(my_filter_reg_coefficients_n93)
         );
  OAI21_X1 my_filter_reg_coefficients_U159 ( .B1(
        my_filter_reg_coefficients_n473), .B2(my_filter_reg_coefficients_n196), 
        .A(my_filter_reg_coefficients_n93), .ZN(
        my_filter_reg_coefficients_n401) );
  NAND2_X1 my_filter_reg_coefficients_U158 ( .A1(b6[6]), .A2(
        my_filter_reg_coefficients_n486), .ZN(my_filter_reg_coefficients_n94)
         );
  OAI21_X1 my_filter_reg_coefficients_U157 ( .B1(
        my_filter_reg_coefficients_n473), .B2(my_filter_reg_coefficients_n195), 
        .A(my_filter_reg_coefficients_n94), .ZN(
        my_filter_reg_coefficients_n402) );
  NAND2_X1 my_filter_reg_coefficients_U156 ( .A1(b6[5]), .A2(
        my_filter_reg_coefficients_n486), .ZN(my_filter_reg_coefficients_n95)
         );
  OAI21_X1 my_filter_reg_coefficients_U155 ( .B1(
        my_filter_reg_coefficients_n473), .B2(my_filter_reg_coefficients_n194), 
        .A(my_filter_reg_coefficients_n95), .ZN(
        my_filter_reg_coefficients_n403) );
  NAND2_X1 my_filter_reg_coefficients_U154 ( .A1(b6[4]), .A2(
        my_filter_reg_coefficients_n486), .ZN(my_filter_reg_coefficients_n96)
         );
  OAI21_X1 my_filter_reg_coefficients_U153 ( .B1(
        my_filter_reg_coefficients_n473), .B2(my_filter_reg_coefficients_n193), 
        .A(my_filter_reg_coefficients_n96), .ZN(
        my_filter_reg_coefficients_n404) );
  NAND2_X1 my_filter_reg_coefficients_U152 ( .A1(b6[3]), .A2(
        my_filter_reg_coefficients_n485), .ZN(my_filter_reg_coefficients_n97)
         );
  OAI21_X1 my_filter_reg_coefficients_U151 ( .B1(
        my_filter_reg_coefficients_n472), .B2(my_filter_reg_coefficients_n192), 
        .A(my_filter_reg_coefficients_n97), .ZN(
        my_filter_reg_coefficients_n405) );
  NAND2_X1 my_filter_reg_coefficients_U150 ( .A1(b6[2]), .A2(
        my_filter_reg_coefficients_n485), .ZN(my_filter_reg_coefficients_n98)
         );
  OAI21_X1 my_filter_reg_coefficients_U149 ( .B1(
        my_filter_reg_coefficients_n472), .B2(my_filter_reg_coefficients_n191), 
        .A(my_filter_reg_coefficients_n98), .ZN(
        my_filter_reg_coefficients_n406) );
  NAND2_X1 my_filter_reg_coefficients_U148 ( .A1(b6[1]), .A2(
        my_filter_reg_coefficients_n485), .ZN(my_filter_reg_coefficients_n99)
         );
  OAI21_X1 my_filter_reg_coefficients_U147 ( .B1(
        my_filter_reg_coefficients_n472), .B2(my_filter_reg_coefficients_n190), 
        .A(my_filter_reg_coefficients_n99), .ZN(
        my_filter_reg_coefficients_n407) );
  NAND2_X1 my_filter_reg_coefficients_U146 ( .A1(b6[0]), .A2(
        my_filter_reg_coefficients_n485), .ZN(my_filter_reg_coefficients_n100)
         );
  OAI21_X1 my_filter_reg_coefficients_U145 ( .B1(
        my_filter_reg_coefficients_n472), .B2(my_filter_reg_coefficients_n189), 
        .A(my_filter_reg_coefficients_n100), .ZN(
        my_filter_reg_coefficients_n408) );
  NAND2_X1 my_filter_reg_coefficients_U144 ( .A1(b7[13]), .A2(
        my_filter_reg_coefficients_n485), .ZN(my_filter_reg_coefficients_n101)
         );
  OAI21_X1 my_filter_reg_coefficients_U143 ( .B1(
        my_filter_reg_coefficients_n472), .B2(my_filter_reg_coefficients_n188), 
        .A(my_filter_reg_coefficients_n101), .ZN(
        my_filter_reg_coefficients_n409) );
  NAND2_X1 my_filter_reg_coefficients_U142 ( .A1(b7[12]), .A2(
        my_filter_reg_coefficients_n485), .ZN(my_filter_reg_coefficients_n102)
         );
  OAI21_X1 my_filter_reg_coefficients_U141 ( .B1(
        my_filter_reg_coefficients_n472), .B2(my_filter_reg_coefficients_n187), 
        .A(my_filter_reg_coefficients_n102), .ZN(
        my_filter_reg_coefficients_n410) );
  NAND2_X1 my_filter_reg_coefficients_U140 ( .A1(b7[11]), .A2(
        my_filter_reg_coefficients_n485), .ZN(my_filter_reg_coefficients_n103)
         );
  OAI21_X1 my_filter_reg_coefficients_U139 ( .B1(
        my_filter_reg_coefficients_n472), .B2(my_filter_reg_coefficients_n186), 
        .A(my_filter_reg_coefficients_n103), .ZN(
        my_filter_reg_coefficients_n411) );
  NAND2_X1 my_filter_reg_coefficients_U138 ( .A1(b7[10]), .A2(
        my_filter_reg_coefficients_n485), .ZN(my_filter_reg_coefficients_n104)
         );
  OAI21_X1 my_filter_reg_coefficients_U137 ( .B1(
        my_filter_reg_coefficients_n472), .B2(my_filter_reg_coefficients_n185), 
        .A(my_filter_reg_coefficients_n104), .ZN(
        my_filter_reg_coefficients_n412) );
  NAND2_X1 my_filter_reg_coefficients_U136 ( .A1(b7[9]), .A2(
        my_filter_reg_coefficients_n485), .ZN(my_filter_reg_coefficients_n105)
         );
  OAI21_X1 my_filter_reg_coefficients_U135 ( .B1(
        my_filter_reg_coefficients_n472), .B2(my_filter_reg_coefficients_n184), 
        .A(my_filter_reg_coefficients_n105), .ZN(
        my_filter_reg_coefficients_n413) );
  NAND2_X1 my_filter_reg_coefficients_U134 ( .A1(b7[8]), .A2(
        my_filter_reg_coefficients_n485), .ZN(my_filter_reg_coefficients_n106)
         );
  OAI21_X1 my_filter_reg_coefficients_U133 ( .B1(
        my_filter_reg_coefficients_n472), .B2(my_filter_reg_coefficients_n183), 
        .A(my_filter_reg_coefficients_n106), .ZN(
        my_filter_reg_coefficients_n414) );
  NAND2_X1 my_filter_reg_coefficients_U132 ( .A1(b7[7]), .A2(
        my_filter_reg_coefficients_n485), .ZN(my_filter_reg_coefficients_n107)
         );
  OAI21_X1 my_filter_reg_coefficients_U131 ( .B1(
        my_filter_reg_coefficients_n472), .B2(my_filter_reg_coefficients_n182), 
        .A(my_filter_reg_coefficients_n107), .ZN(
        my_filter_reg_coefficients_n415) );
  NAND2_X1 my_filter_reg_coefficients_U130 ( .A1(b7[6]), .A2(
        my_filter_reg_coefficients_n485), .ZN(my_filter_reg_coefficients_n108)
         );
  OAI21_X1 my_filter_reg_coefficients_U129 ( .B1(
        my_filter_reg_coefficients_n472), .B2(my_filter_reg_coefficients_n181), 
        .A(my_filter_reg_coefficients_n108), .ZN(
        my_filter_reg_coefficients_n416) );
  NAND2_X1 my_filter_reg_coefficients_U128 ( .A1(b7[5]), .A2(
        my_filter_reg_coefficients_n484), .ZN(my_filter_reg_coefficients_n109)
         );
  OAI21_X1 my_filter_reg_coefficients_U127 ( .B1(
        my_filter_reg_coefficients_n471), .B2(my_filter_reg_coefficients_n180), 
        .A(my_filter_reg_coefficients_n109), .ZN(
        my_filter_reg_coefficients_n417) );
  NAND2_X1 my_filter_reg_coefficients_U126 ( .A1(b7[4]), .A2(
        my_filter_reg_coefficients_n484), .ZN(my_filter_reg_coefficients_n110)
         );
  OAI21_X1 my_filter_reg_coefficients_U125 ( .B1(
        my_filter_reg_coefficients_n471), .B2(my_filter_reg_coefficients_n179), 
        .A(my_filter_reg_coefficients_n110), .ZN(
        my_filter_reg_coefficients_n418) );
  NAND2_X1 my_filter_reg_coefficients_U124 ( .A1(b7[3]), .A2(
        my_filter_reg_coefficients_n484), .ZN(my_filter_reg_coefficients_n111)
         );
  OAI21_X1 my_filter_reg_coefficients_U123 ( .B1(
        my_filter_reg_coefficients_n471), .B2(my_filter_reg_coefficients_n178), 
        .A(my_filter_reg_coefficients_n111), .ZN(
        my_filter_reg_coefficients_n419) );
  NAND2_X1 my_filter_reg_coefficients_U122 ( .A1(b7[2]), .A2(
        my_filter_reg_coefficients_n484), .ZN(my_filter_reg_coefficients_n112)
         );
  OAI21_X1 my_filter_reg_coefficients_U121 ( .B1(
        my_filter_reg_coefficients_n471), .B2(my_filter_reg_coefficients_n177), 
        .A(my_filter_reg_coefficients_n112), .ZN(
        my_filter_reg_coefficients_n420) );
  NAND2_X1 my_filter_reg_coefficients_U120 ( .A1(b7[1]), .A2(
        my_filter_reg_coefficients_n484), .ZN(my_filter_reg_coefficients_n113)
         );
  OAI21_X1 my_filter_reg_coefficients_U119 ( .B1(
        my_filter_reg_coefficients_n471), .B2(my_filter_reg_coefficients_n176), 
        .A(my_filter_reg_coefficients_n113), .ZN(
        my_filter_reg_coefficients_n421) );
  NAND2_X1 my_filter_reg_coefficients_U118 ( .A1(b7[0]), .A2(
        my_filter_reg_coefficients_n484), .ZN(my_filter_reg_coefficients_n114)
         );
  OAI21_X1 my_filter_reg_coefficients_U117 ( .B1(
        my_filter_reg_coefficients_n471), .B2(my_filter_reg_coefficients_n175), 
        .A(my_filter_reg_coefficients_n114), .ZN(
        my_filter_reg_coefficients_n422) );
  NAND2_X1 my_filter_reg_coefficients_U116 ( .A1(b8[13]), .A2(
        my_filter_reg_coefficients_n484), .ZN(my_filter_reg_coefficients_n115)
         );
  OAI21_X1 my_filter_reg_coefficients_U115 ( .B1(
        my_filter_reg_coefficients_n471), .B2(my_filter_reg_coefficients_n174), 
        .A(my_filter_reg_coefficients_n115), .ZN(
        my_filter_reg_coefficients_n423) );
  NAND2_X1 my_filter_reg_coefficients_U114 ( .A1(b8[12]), .A2(
        my_filter_reg_coefficients_n484), .ZN(my_filter_reg_coefficients_n116)
         );
  OAI21_X1 my_filter_reg_coefficients_U113 ( .B1(
        my_filter_reg_coefficients_n471), .B2(my_filter_reg_coefficients_n173), 
        .A(my_filter_reg_coefficients_n116), .ZN(
        my_filter_reg_coefficients_n424) );
  NAND2_X1 my_filter_reg_coefficients_U112 ( .A1(b8[11]), .A2(
        my_filter_reg_coefficients_n484), .ZN(my_filter_reg_coefficients_n117)
         );
  OAI21_X1 my_filter_reg_coefficients_U111 ( .B1(
        my_filter_reg_coefficients_n471), .B2(my_filter_reg_coefficients_n172), 
        .A(my_filter_reg_coefficients_n117), .ZN(
        my_filter_reg_coefficients_n425) );
  NAND2_X1 my_filter_reg_coefficients_U110 ( .A1(b8[10]), .A2(
        my_filter_reg_coefficients_n484), .ZN(my_filter_reg_coefficients_n118)
         );
  OAI21_X1 my_filter_reg_coefficients_U109 ( .B1(
        my_filter_reg_coefficients_n471), .B2(my_filter_reg_coefficients_n171), 
        .A(my_filter_reg_coefficients_n118), .ZN(
        my_filter_reg_coefficients_n426) );
  NAND2_X1 my_filter_reg_coefficients_U108 ( .A1(b8[9]), .A2(
        my_filter_reg_coefficients_n484), .ZN(my_filter_reg_coefficients_n119)
         );
  OAI21_X1 my_filter_reg_coefficients_U107 ( .B1(
        my_filter_reg_coefficients_n471), .B2(my_filter_reg_coefficients_n170), 
        .A(my_filter_reg_coefficients_n119), .ZN(
        my_filter_reg_coefficients_n427) );
  NAND2_X1 my_filter_reg_coefficients_U106 ( .A1(b8[8]), .A2(
        my_filter_reg_coefficients_n484), .ZN(my_filter_reg_coefficients_n120)
         );
  OAI21_X1 my_filter_reg_coefficients_U105 ( .B1(
        my_filter_reg_coefficients_n471), .B2(my_filter_reg_coefficients_n169), 
        .A(my_filter_reg_coefficients_n120), .ZN(
        my_filter_reg_coefficients_n428) );
  NAND2_X1 my_filter_reg_coefficients_U104 ( .A1(b8[7]), .A2(
        my_filter_reg_coefficients_n483), .ZN(my_filter_reg_coefficients_n121)
         );
  OAI21_X1 my_filter_reg_coefficients_U103 ( .B1(
        my_filter_reg_coefficients_n470), .B2(my_filter_reg_coefficients_n168), 
        .A(my_filter_reg_coefficients_n121), .ZN(
        my_filter_reg_coefficients_n429) );
  NAND2_X1 my_filter_reg_coefficients_U102 ( .A1(b8[6]), .A2(
        my_filter_reg_coefficients_n483), .ZN(my_filter_reg_coefficients_n122)
         );
  OAI21_X1 my_filter_reg_coefficients_U101 ( .B1(
        my_filter_reg_coefficients_n470), .B2(my_filter_reg_coefficients_n167), 
        .A(my_filter_reg_coefficients_n122), .ZN(
        my_filter_reg_coefficients_n430) );
  NAND2_X1 my_filter_reg_coefficients_U100 ( .A1(b8[5]), .A2(
        my_filter_reg_coefficients_n483), .ZN(my_filter_reg_coefficients_n123)
         );
  OAI21_X1 my_filter_reg_coefficients_U99 ( .B1(
        my_filter_reg_coefficients_n470), .B2(my_filter_reg_coefficients_n310), 
        .A(my_filter_reg_coefficients_n123), .ZN(
        my_filter_reg_coefficients_n431) );
  NAND2_X1 my_filter_reg_coefficients_U98 ( .A1(b8[4]), .A2(
        my_filter_reg_coefficients_n483), .ZN(my_filter_reg_coefficients_n124)
         );
  OAI21_X1 my_filter_reg_coefficients_U97 ( .B1(
        my_filter_reg_coefficients_n470), .B2(my_filter_reg_coefficients_n309), 
        .A(my_filter_reg_coefficients_n124), .ZN(
        my_filter_reg_coefficients_n432) );
  NAND2_X1 my_filter_reg_coefficients_U96 ( .A1(b8[3]), .A2(
        my_filter_reg_coefficients_n483), .ZN(my_filter_reg_coefficients_n125)
         );
  OAI21_X1 my_filter_reg_coefficients_U95 ( .B1(
        my_filter_reg_coefficients_n470), .B2(my_filter_reg_coefficients_n308), 
        .A(my_filter_reg_coefficients_n125), .ZN(
        my_filter_reg_coefficients_n433) );
  NAND2_X1 my_filter_reg_coefficients_U94 ( .A1(b8[2]), .A2(
        my_filter_reg_coefficients_n483), .ZN(my_filter_reg_coefficients_n126)
         );
  OAI21_X1 my_filter_reg_coefficients_U93 ( .B1(
        my_filter_reg_coefficients_n470), .B2(my_filter_reg_coefficients_n307), 
        .A(my_filter_reg_coefficients_n126), .ZN(
        my_filter_reg_coefficients_n434) );
  NAND2_X1 my_filter_reg_coefficients_U92 ( .A1(b8[1]), .A2(
        my_filter_reg_coefficients_n483), .ZN(my_filter_reg_coefficients_n127)
         );
  OAI21_X1 my_filter_reg_coefficients_U91 ( .B1(
        my_filter_reg_coefficients_n470), .B2(my_filter_reg_coefficients_n306), 
        .A(my_filter_reg_coefficients_n127), .ZN(
        my_filter_reg_coefficients_n435) );
  NAND2_X1 my_filter_reg_coefficients_U90 ( .A1(b8[0]), .A2(
        my_filter_reg_coefficients_n483), .ZN(my_filter_reg_coefficients_n128)
         );
  OAI21_X1 my_filter_reg_coefficients_U89 ( .B1(
        my_filter_reg_coefficients_n470), .B2(my_filter_reg_coefficients_n290), 
        .A(my_filter_reg_coefficients_n128), .ZN(
        my_filter_reg_coefficients_n436) );
  NAND2_X1 my_filter_reg_coefficients_U88 ( .A1(b9[13]), .A2(
        my_filter_reg_coefficients_n483), .ZN(my_filter_reg_coefficients_n129)
         );
  OAI21_X1 my_filter_reg_coefficients_U87 ( .B1(
        my_filter_reg_coefficients_n470), .B2(my_filter_reg_coefficients_n288), 
        .A(my_filter_reg_coefficients_n129), .ZN(
        my_filter_reg_coefficients_n437) );
  NAND2_X1 my_filter_reg_coefficients_U86 ( .A1(b9[12]), .A2(
        my_filter_reg_coefficients_n483), .ZN(my_filter_reg_coefficients_n130)
         );
  OAI21_X1 my_filter_reg_coefficients_U85 ( .B1(
        my_filter_reg_coefficients_n470), .B2(my_filter_reg_coefficients_n305), 
        .A(my_filter_reg_coefficients_n130), .ZN(
        my_filter_reg_coefficients_n438) );
  NAND2_X1 my_filter_reg_coefficients_U84 ( .A1(b9[11]), .A2(
        my_filter_reg_coefficients_n483), .ZN(my_filter_reg_coefficients_n131)
         );
  OAI21_X1 my_filter_reg_coefficients_U83 ( .B1(
        my_filter_reg_coefficients_n470), .B2(my_filter_reg_coefficients_n304), 
        .A(my_filter_reg_coefficients_n131), .ZN(
        my_filter_reg_coefficients_n439) );
  NAND2_X1 my_filter_reg_coefficients_U82 ( .A1(b9[10]), .A2(
        my_filter_reg_coefficients_n483), .ZN(my_filter_reg_coefficients_n132)
         );
  OAI21_X1 my_filter_reg_coefficients_U81 ( .B1(
        my_filter_reg_coefficients_n470), .B2(my_filter_reg_coefficients_n303), 
        .A(my_filter_reg_coefficients_n132), .ZN(
        my_filter_reg_coefficients_n440) );
  NAND2_X1 my_filter_reg_coefficients_U80 ( .A1(b9[9]), .A2(
        my_filter_reg_coefficients_n482), .ZN(my_filter_reg_coefficients_n133)
         );
  OAI21_X1 my_filter_reg_coefficients_U79 ( .B1(
        my_filter_reg_coefficients_n469), .B2(my_filter_reg_coefficients_n302), 
        .A(my_filter_reg_coefficients_n133), .ZN(
        my_filter_reg_coefficients_n441) );
  NAND2_X1 my_filter_reg_coefficients_U78 ( .A1(b9[8]), .A2(
        my_filter_reg_coefficients_n482), .ZN(my_filter_reg_coefficients_n134)
         );
  OAI21_X1 my_filter_reg_coefficients_U77 ( .B1(
        my_filter_reg_coefficients_n469), .B2(my_filter_reg_coefficients_n301), 
        .A(my_filter_reg_coefficients_n134), .ZN(
        my_filter_reg_coefficients_n442) );
  NAND2_X1 my_filter_reg_coefficients_U76 ( .A1(b9[7]), .A2(
        my_filter_reg_coefficients_n482), .ZN(my_filter_reg_coefficients_n135)
         );
  OAI21_X1 my_filter_reg_coefficients_U75 ( .B1(
        my_filter_reg_coefficients_n469), .B2(my_filter_reg_coefficients_n300), 
        .A(my_filter_reg_coefficients_n135), .ZN(
        my_filter_reg_coefficients_n443) );
  NAND2_X1 my_filter_reg_coefficients_U74 ( .A1(b9[6]), .A2(
        my_filter_reg_coefficients_n482), .ZN(my_filter_reg_coefficients_n136)
         );
  OAI21_X1 my_filter_reg_coefficients_U73 ( .B1(
        my_filter_reg_coefficients_n469), .B2(my_filter_reg_coefficients_n299), 
        .A(my_filter_reg_coefficients_n136), .ZN(
        my_filter_reg_coefficients_n444) );
  NAND2_X1 my_filter_reg_coefficients_U72 ( .A1(b9[5]), .A2(
        my_filter_reg_coefficients_n482), .ZN(my_filter_reg_coefficients_n137)
         );
  OAI21_X1 my_filter_reg_coefficients_U71 ( .B1(
        my_filter_reg_coefficients_n469), .B2(my_filter_reg_coefficients_n298), 
        .A(my_filter_reg_coefficients_n137), .ZN(
        my_filter_reg_coefficients_n445) );
  NAND2_X1 my_filter_reg_coefficients_U70 ( .A1(b9[4]), .A2(
        my_filter_reg_coefficients_n482), .ZN(my_filter_reg_coefficients_n138)
         );
  OAI21_X1 my_filter_reg_coefficients_U69 ( .B1(
        my_filter_reg_coefficients_n469), .B2(my_filter_reg_coefficients_n297), 
        .A(my_filter_reg_coefficients_n138), .ZN(
        my_filter_reg_coefficients_n446) );
  NAND2_X1 my_filter_reg_coefficients_U68 ( .A1(b9[3]), .A2(
        my_filter_reg_coefficients_n482), .ZN(my_filter_reg_coefficients_n139)
         );
  OAI21_X1 my_filter_reg_coefficients_U67 ( .B1(
        my_filter_reg_coefficients_n469), .B2(my_filter_reg_coefficients_n296), 
        .A(my_filter_reg_coefficients_n139), .ZN(
        my_filter_reg_coefficients_n447) );
  NAND2_X1 my_filter_reg_coefficients_U66 ( .A1(b9[2]), .A2(
        my_filter_reg_coefficients_n482), .ZN(my_filter_reg_coefficients_n140)
         );
  OAI21_X1 my_filter_reg_coefficients_U65 ( .B1(
        my_filter_reg_coefficients_n469), .B2(my_filter_reg_coefficients_n295), 
        .A(my_filter_reg_coefficients_n140), .ZN(
        my_filter_reg_coefficients_n448) );
  NAND2_X1 my_filter_reg_coefficients_U64 ( .A1(b9[1]), .A2(
        my_filter_reg_coefficients_n482), .ZN(my_filter_reg_coefficients_n141)
         );
  OAI21_X1 my_filter_reg_coefficients_U63 ( .B1(
        my_filter_reg_coefficients_n469), .B2(my_filter_reg_coefficients_n294), 
        .A(my_filter_reg_coefficients_n141), .ZN(
        my_filter_reg_coefficients_n449) );
  NAND2_X1 my_filter_reg_coefficients_U62 ( .A1(b9[0]), .A2(
        my_filter_reg_coefficients_n482), .ZN(my_filter_reg_coefficients_n142)
         );
  OAI21_X1 my_filter_reg_coefficients_U61 ( .B1(
        my_filter_reg_coefficients_n469), .B2(my_filter_reg_coefficients_n289), 
        .A(my_filter_reg_coefficients_n142), .ZN(
        my_filter_reg_coefficients_n450) );
  NAND2_X1 my_filter_reg_coefficients_U60 ( .A1(b10[13]), .A2(
        my_filter_reg_coefficients_n482), .ZN(my_filter_reg_coefficients_n143)
         );
  OAI21_X1 my_filter_reg_coefficients_U59 ( .B1(
        my_filter_reg_coefficients_n469), .B2(my_filter_reg_coefficients_n287), 
        .A(my_filter_reg_coefficients_n143), .ZN(
        my_filter_reg_coefficients_n451) );
  NAND2_X1 my_filter_reg_coefficients_U58 ( .A1(b10[12]), .A2(
        my_filter_reg_coefficients_n482), .ZN(my_filter_reg_coefficients_n144)
         );
  OAI21_X1 my_filter_reg_coefficients_U57 ( .B1(
        my_filter_reg_coefficients_n469), .B2(my_filter_reg_coefficients_n293), 
        .A(my_filter_reg_coefficients_n144), .ZN(
        my_filter_reg_coefficients_n452) );
  NAND2_X1 my_filter_reg_coefficients_U56 ( .A1(b10[11]), .A2(
        my_filter_reg_coefficients_n481), .ZN(my_filter_reg_coefficients_n145)
         );
  OAI21_X1 my_filter_reg_coefficients_U55 ( .B1(
        my_filter_reg_coefficients_n468), .B2(my_filter_reg_coefficients_n292), 
        .A(my_filter_reg_coefficients_n145), .ZN(
        my_filter_reg_coefficients_n453) );
  NAND2_X1 my_filter_reg_coefficients_U54 ( .A1(b10[10]), .A2(
        my_filter_reg_coefficients_n481), .ZN(my_filter_reg_coefficients_n146)
         );
  OAI21_X1 my_filter_reg_coefficients_U53 ( .B1(
        my_filter_reg_coefficients_n468), .B2(my_filter_reg_coefficients_n291), 
        .A(my_filter_reg_coefficients_n146), .ZN(
        my_filter_reg_coefficients_n454) );
  NAND2_X1 my_filter_reg_coefficients_U52 ( .A1(b10[9]), .A2(
        my_filter_reg_coefficients_n481), .ZN(my_filter_reg_coefficients_n147)
         );
  OAI21_X1 my_filter_reg_coefficients_U51 ( .B1(
        my_filter_reg_coefficients_n468), .B2(my_filter_reg_coefficients_n166), 
        .A(my_filter_reg_coefficients_n147), .ZN(
        my_filter_reg_coefficients_n455) );
  NAND2_X1 my_filter_reg_coefficients_U50 ( .A1(b10[8]), .A2(
        my_filter_reg_coefficients_n481), .ZN(my_filter_reg_coefficients_n148)
         );
  OAI21_X1 my_filter_reg_coefficients_U49 ( .B1(
        my_filter_reg_coefficients_n468), .B2(my_filter_reg_coefficients_n165), 
        .A(my_filter_reg_coefficients_n148), .ZN(
        my_filter_reg_coefficients_n456) );
  NAND2_X1 my_filter_reg_coefficients_U48 ( .A1(b10[7]), .A2(
        my_filter_reg_coefficients_n481), .ZN(my_filter_reg_coefficients_n149)
         );
  OAI21_X1 my_filter_reg_coefficients_U47 ( .B1(
        my_filter_reg_coefficients_n468), .B2(my_filter_reg_coefficients_n164), 
        .A(my_filter_reg_coefficients_n149), .ZN(
        my_filter_reg_coefficients_n457) );
  NAND2_X1 my_filter_reg_coefficients_U46 ( .A1(b10[6]), .A2(
        my_filter_reg_coefficients_n481), .ZN(my_filter_reg_coefficients_n150)
         );
  OAI21_X1 my_filter_reg_coefficients_U45 ( .B1(
        my_filter_reg_coefficients_n468), .B2(my_filter_reg_coefficients_n163), 
        .A(my_filter_reg_coefficients_n150), .ZN(
        my_filter_reg_coefficients_n458) );
  NAND2_X1 my_filter_reg_coefficients_U44 ( .A1(b10[5]), .A2(
        my_filter_reg_coefficients_n481), .ZN(my_filter_reg_coefficients_n151)
         );
  OAI21_X1 my_filter_reg_coefficients_U43 ( .B1(
        my_filter_reg_coefficients_n468), .B2(my_filter_reg_coefficients_n162), 
        .A(my_filter_reg_coefficients_n151), .ZN(
        my_filter_reg_coefficients_n459) );
  NAND2_X1 my_filter_reg_coefficients_U42 ( .A1(b10[4]), .A2(
        my_filter_reg_coefficients_n481), .ZN(my_filter_reg_coefficients_n152)
         );
  OAI21_X1 my_filter_reg_coefficients_U41 ( .B1(
        my_filter_reg_coefficients_n468), .B2(my_filter_reg_coefficients_n161), 
        .A(my_filter_reg_coefficients_n152), .ZN(
        my_filter_reg_coefficients_n460) );
  NAND2_X1 my_filter_reg_coefficients_U40 ( .A1(b10[3]), .A2(
        my_filter_reg_coefficients_n481), .ZN(my_filter_reg_coefficients_n153)
         );
  OAI21_X1 my_filter_reg_coefficients_U39 ( .B1(
        my_filter_reg_coefficients_n468), .B2(my_filter_reg_coefficients_n160), 
        .A(my_filter_reg_coefficients_n153), .ZN(
        my_filter_reg_coefficients_n461) );
  NAND2_X1 my_filter_reg_coefficients_U38 ( .A1(b10[2]), .A2(
        my_filter_reg_coefficients_n481), .ZN(my_filter_reg_coefficients_n154)
         );
  OAI21_X1 my_filter_reg_coefficients_U37 ( .B1(
        my_filter_reg_coefficients_n468), .B2(my_filter_reg_coefficients_n159), 
        .A(my_filter_reg_coefficients_n154), .ZN(
        my_filter_reg_coefficients_n462) );
  NAND2_X1 my_filter_reg_coefficients_U36 ( .A1(b10[1]), .A2(
        my_filter_reg_coefficients_n481), .ZN(my_filter_reg_coefficients_n155)
         );
  OAI21_X1 my_filter_reg_coefficients_U35 ( .B1(
        my_filter_reg_coefficients_n468), .B2(my_filter_reg_coefficients_n158), 
        .A(my_filter_reg_coefficients_n155), .ZN(
        my_filter_reg_coefficients_n463) );
  NAND2_X1 my_filter_reg_coefficients_U34 ( .A1(b10[0]), .A2(
        my_filter_reg_coefficients_n481), .ZN(my_filter_reg_coefficients_n156)
         );
  OAI21_X1 my_filter_reg_coefficients_U33 ( .B1(
        my_filter_reg_coefficients_n468), .B2(my_filter_reg_coefficients_n157), 
        .A(my_filter_reg_coefficients_n156), .ZN(
        my_filter_reg_coefficients_n464) );
  INV_X1 my_filter_reg_coefficients_U32 ( .A(my_filter_reg_coefficients_n493), 
        .ZN(my_filter_reg_coefficients_n492) );
  INV_X1 my_filter_reg_coefficients_U31 ( .A(my_filter_reg_coefficients_n493), 
        .ZN(my_filter_reg_coefficients_n491) );
  INV_X1 my_filter_reg_coefficients_U30 ( .A(my_filter_reg_coefficients_n493), 
        .ZN(my_filter_reg_coefficients_n490) );
  INV_X1 my_filter_reg_coefficients_U29 ( .A(my_filter_reg_coefficients_n493), 
        .ZN(my_filter_reg_coefficients_n489) );
  INV_X1 my_filter_reg_coefficients_U28 ( .A(my_filter_reg_coefficients_n493), 
        .ZN(my_filter_reg_coefficients_n488) );
  INV_X1 my_filter_reg_coefficients_U27 ( .A(my_filter_reg_coefficients_n493), 
        .ZN(my_filter_reg_coefficients_n487) );
  INV_X1 my_filter_reg_coefficients_U26 ( .A(my_filter_reg_coefficients_n493), 
        .ZN(my_filter_reg_coefficients_n486) );
  INV_X1 my_filter_reg_coefficients_U25 ( .A(my_filter_reg_coefficients_n493), 
        .ZN(my_filter_reg_coefficients_n485) );
  INV_X1 my_filter_reg_coefficients_U24 ( .A(my_filter_reg_coefficients_n493), 
        .ZN(my_filter_reg_coefficients_n484) );
  INV_X1 my_filter_reg_coefficients_U23 ( .A(my_filter_reg_coefficients_n493), 
        .ZN(my_filter_reg_coefficients_n483) );
  INV_X1 my_filter_reg_coefficients_U22 ( .A(my_filter_reg_coefficients_n493), 
        .ZN(my_filter_reg_coefficients_n482) );
  INV_X1 my_filter_reg_coefficients_U21 ( .A(my_filter_reg_coefficients_n493), 
        .ZN(my_filter_reg_coefficients_n481) );
  NAND2_X1 my_filter_reg_coefficients_U20 ( .A1(
        my_filter_reg_coefficients_n497), .A2(my_filter_reg_coefficients_n493), 
        .ZN(my_filter_reg_coefficients_n2) );
  BUF_X1 my_filter_reg_coefficients_U19 ( .A(my_filter_reg_coefficients_n2), 
        .Z(my_filter_reg_coefficients_n467) );
  BUF_X1 my_filter_reg_coefficients_U18 ( .A(my_filter_reg_coefficients_n2), 
        .Z(my_filter_reg_coefficients_n466) );
  BUF_X1 my_filter_reg_coefficients_U17 ( .A(my_filter_reg_coefficients_n2), 
        .Z(my_filter_reg_coefficients_n465) );
  BUF_X1 my_filter_reg_coefficients_U16 ( .A(my_filter_reg_coefficients_n494), 
        .Z(my_filter_reg_coefficients_n497) );
  BUF_X1 my_filter_reg_coefficients_U15 ( .A(my_filter_reg_coefficients_n467), 
        .Z(my_filter_reg_coefficients_n480) );
  BUF_X1 my_filter_reg_coefficients_U14 ( .A(my_filter_reg_coefficients_n467), 
        .Z(my_filter_reg_coefficients_n479) );
  BUF_X1 my_filter_reg_coefficients_U13 ( .A(my_filter_reg_coefficients_n467), 
        .Z(my_filter_reg_coefficients_n478) );
  BUF_X1 my_filter_reg_coefficients_U12 ( .A(my_filter_reg_coefficients_n466), 
        .Z(my_filter_reg_coefficients_n477) );
  BUF_X1 my_filter_reg_coefficients_U11 ( .A(my_filter_reg_coefficients_n466), 
        .Z(my_filter_reg_coefficients_n476) );
  BUF_X1 my_filter_reg_coefficients_U10 ( .A(my_filter_reg_coefficients_n466), 
        .Z(my_filter_reg_coefficients_n475) );
  BUF_X1 my_filter_reg_coefficients_U9 ( .A(my_filter_reg_coefficients_n466), 
        .Z(my_filter_reg_coefficients_n474) );
  BUF_X1 my_filter_reg_coefficients_U8 ( .A(my_filter_reg_coefficients_n466), 
        .Z(my_filter_reg_coefficients_n473) );
  BUF_X1 my_filter_reg_coefficients_U7 ( .A(my_filter_reg_coefficients_n465), 
        .Z(my_filter_reg_coefficients_n472) );
  BUF_X1 my_filter_reg_coefficients_U6 ( .A(my_filter_reg_coefficients_n465), 
        .Z(my_filter_reg_coefficients_n471) );
  BUF_X1 my_filter_reg_coefficients_U5 ( .A(my_filter_reg_coefficients_n465), 
        .Z(my_filter_reg_coefficients_n470) );
  BUF_X1 my_filter_reg_coefficients_U4 ( .A(my_filter_reg_coefficients_n465), 
        .Z(my_filter_reg_coefficients_n469) );
  BUF_X1 my_filter_reg_coefficients_U3 ( .A(my_filter_reg_coefficients_n465), 
        .Z(my_filter_reg_coefficients_n468) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_10__0_ ( .D(
        my_filter_reg_coefficients_n464), .CK(clk), .RN(
        my_filter_reg_coefficients_n503), .Q(my_filter_q_reg_coeff[0]), .QN(
        my_filter_reg_coefficients_n157) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_10__1_ ( .D(
        my_filter_reg_coefficients_n463), .CK(clk), .RN(
        my_filter_reg_coefficients_n503), .Q(my_filter_q_reg_coeff[1]), .QN(
        my_filter_reg_coefficients_n158) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_10__2_ ( .D(
        my_filter_reg_coefficients_n462), .CK(clk), .RN(
        my_filter_reg_coefficients_n503), .Q(my_filter_q_reg_coeff[2]), .QN(
        my_filter_reg_coefficients_n159) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_10__3_ ( .D(
        my_filter_reg_coefficients_n461), .CK(clk), .RN(
        my_filter_reg_coefficients_n503), .Q(my_filter_q_reg_coeff[3]), .QN(
        my_filter_reg_coefficients_n160) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_10__4_ ( .D(
        my_filter_reg_coefficients_n460), .CK(clk), .RN(
        my_filter_reg_coefficients_n503), .Q(my_filter_q_reg_coeff[4]), .QN(
        my_filter_reg_coefficients_n161) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_10__5_ ( .D(
        my_filter_reg_coefficients_n459), .CK(clk), .RN(
        my_filter_reg_coefficients_n503), .Q(my_filter_q_reg_coeff[5]), .QN(
        my_filter_reg_coefficients_n162) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_10__6_ ( .D(
        my_filter_reg_coefficients_n458), .CK(clk), .RN(
        my_filter_reg_coefficients_n503), .Q(my_filter_q_reg_coeff[6]), .QN(
        my_filter_reg_coefficients_n163) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_10__7_ ( .D(
        my_filter_reg_coefficients_n457), .CK(clk), .RN(
        my_filter_reg_coefficients_n503), .Q(my_filter_q_reg_coeff[7]), .QN(
        my_filter_reg_coefficients_n164) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_10__8_ ( .D(
        my_filter_reg_coefficients_n456), .CK(clk), .RN(
        my_filter_reg_coefficients_n503), .Q(my_filter_q_reg_coeff[8]), .QN(
        my_filter_reg_coefficients_n165) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_10__9_ ( .D(
        my_filter_reg_coefficients_n455), .CK(clk), .RN(
        my_filter_reg_coefficients_n503), .Q(my_filter_q_reg_coeff[9]), .QN(
        my_filter_reg_coefficients_n166) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_10__10_ ( .D(
        my_filter_reg_coefficients_n454), .CK(clk), .RN(
        my_filter_reg_coefficients_n503), .Q(my_filter_q_reg_coeff[10]), .QN(
        my_filter_reg_coefficients_n291) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_10__11_ ( .D(
        my_filter_reg_coefficients_n453), .CK(clk), .RN(
        my_filter_reg_coefficients_n503), .Q(my_filter_q_reg_coeff[11]), .QN(
        my_filter_reg_coefficients_n292) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_10__12_ ( .D(
        my_filter_reg_coefficients_n452), .CK(clk), .RN(
        my_filter_reg_coefficients_n503), .Q(my_filter_q_reg_coeff[12]), .QN(
        my_filter_reg_coefficients_n293) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_10__13_ ( .D(
        my_filter_reg_coefficients_n451), .CK(clk), .RN(
        my_filter_reg_coefficients_n503), .Q(my_filter_q_reg_coeff[13]), .QN(
        my_filter_reg_coefficients_n287) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_9__0_ ( .D(
        my_filter_reg_coefficients_n450), .CK(clk), .RN(
        my_filter_reg_coefficients_n502), .Q(my_filter_q_reg_coeff[14]), .QN(
        my_filter_reg_coefficients_n289) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_9__1_ ( .D(
        my_filter_reg_coefficients_n449), .CK(clk), .RN(
        my_filter_reg_coefficients_n502), .Q(my_filter_q_reg_coeff[15]), .QN(
        my_filter_reg_coefficients_n294) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_9__2_ ( .D(
        my_filter_reg_coefficients_n448), .CK(clk), .RN(
        my_filter_reg_coefficients_n502), .Q(my_filter_q_reg_coeff[16]), .QN(
        my_filter_reg_coefficients_n295) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_9__3_ ( .D(
        my_filter_reg_coefficients_n447), .CK(clk), .RN(
        my_filter_reg_coefficients_n502), .Q(my_filter_q_reg_coeff[17]), .QN(
        my_filter_reg_coefficients_n296) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_9__4_ ( .D(
        my_filter_reg_coefficients_n446), .CK(clk), .RN(
        my_filter_reg_coefficients_n502), .Q(my_filter_q_reg_coeff[18]), .QN(
        my_filter_reg_coefficients_n297) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_9__5_ ( .D(
        my_filter_reg_coefficients_n445), .CK(clk), .RN(
        my_filter_reg_coefficients_n502), .Q(my_filter_q_reg_coeff[19]), .QN(
        my_filter_reg_coefficients_n298) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_9__6_ ( .D(
        my_filter_reg_coefficients_n444), .CK(clk), .RN(
        my_filter_reg_coefficients_n502), .Q(my_filter_q_reg_coeff[20]), .QN(
        my_filter_reg_coefficients_n299) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_9__7_ ( .D(
        my_filter_reg_coefficients_n443), .CK(clk), .RN(
        my_filter_reg_coefficients_n502), .Q(my_filter_q_reg_coeff[21]), .QN(
        my_filter_reg_coefficients_n300) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_9__8_ ( .D(
        my_filter_reg_coefficients_n442), .CK(clk), .RN(
        my_filter_reg_coefficients_n502), .Q(my_filter_q_reg_coeff[22]), .QN(
        my_filter_reg_coefficients_n301) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_9__9_ ( .D(
        my_filter_reg_coefficients_n441), .CK(clk), .RN(
        my_filter_reg_coefficients_n502), .Q(my_filter_q_reg_coeff[23]), .QN(
        my_filter_reg_coefficients_n302) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_9__10_ ( .D(
        my_filter_reg_coefficients_n440), .CK(clk), .RN(
        my_filter_reg_coefficients_n502), .Q(my_filter_q_reg_coeff[24]), .QN(
        my_filter_reg_coefficients_n303) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_9__11_ ( .D(
        my_filter_reg_coefficients_n439), .CK(clk), .RN(
        my_filter_reg_coefficients_n502), .Q(my_filter_q_reg_coeff[25]), .QN(
        my_filter_reg_coefficients_n304) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_9__12_ ( .D(
        my_filter_reg_coefficients_n438), .CK(clk), .RN(
        my_filter_reg_coefficients_n502), .Q(my_filter_q_reg_coeff[26]), .QN(
        my_filter_reg_coefficients_n305) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_9__13_ ( .D(
        my_filter_reg_coefficients_n437), .CK(clk), .RN(
        my_filter_reg_coefficients_n502), .Q(my_filter_q_reg_coeff[27]), .QN(
        my_filter_reg_coefficients_n288) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_8__0_ ( .D(
        my_filter_reg_coefficients_n436), .CK(clk), .RN(
        my_filter_reg_coefficients_n501), .Q(my_filter_q_reg_coeff[28]), .QN(
        my_filter_reg_coefficients_n290) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_8__1_ ( .D(
        my_filter_reg_coefficients_n435), .CK(clk), .RN(
        my_filter_reg_coefficients_n501), .Q(my_filter_q_reg_coeff[29]), .QN(
        my_filter_reg_coefficients_n306) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_8__2_ ( .D(
        my_filter_reg_coefficients_n434), .CK(clk), .RN(
        my_filter_reg_coefficients_n502), .Q(my_filter_q_reg_coeff[30]), .QN(
        my_filter_reg_coefficients_n307) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_8__3_ ( .D(
        my_filter_reg_coefficients_n433), .CK(clk), .RN(
        my_filter_reg_coefficients_n502), .Q(my_filter_q_reg_coeff[31]), .QN(
        my_filter_reg_coefficients_n308) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_8__4_ ( .D(
        my_filter_reg_coefficients_n432), .CK(clk), .RN(
        my_filter_reg_coefficients_n502), .Q(my_filter_q_reg_coeff[32]), .QN(
        my_filter_reg_coefficients_n309) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_8__5_ ( .D(
        my_filter_reg_coefficients_n431), .CK(clk), .RN(
        my_filter_reg_coefficients_n502), .Q(my_filter_q_reg_coeff[33]), .QN(
        my_filter_reg_coefficients_n310) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_8__6_ ( .D(
        my_filter_reg_coefficients_n430), .CK(clk), .RN(
        my_filter_reg_coefficients_n501), .Q(my_filter_q_reg_coeff[34]), .QN(
        my_filter_reg_coefficients_n167) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_8__7_ ( .D(
        my_filter_reg_coefficients_n429), .CK(clk), .RN(
        my_filter_reg_coefficients_n501), .Q(my_filter_q_reg_coeff[35]), .QN(
        my_filter_reg_coefficients_n168) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_8__8_ ( .D(
        my_filter_reg_coefficients_n428), .CK(clk), .RN(
        my_filter_reg_coefficients_n501), .Q(my_filter_q_reg_coeff[36]), .QN(
        my_filter_reg_coefficients_n169) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_8__9_ ( .D(
        my_filter_reg_coefficients_n427), .CK(clk), .RN(
        my_filter_reg_coefficients_n501), .Q(my_filter_q_reg_coeff[37]), .QN(
        my_filter_reg_coefficients_n170) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_8__10_ ( .D(
        my_filter_reg_coefficients_n426), .CK(clk), .RN(
        my_filter_reg_coefficients_n501), .Q(my_filter_q_reg_coeff[38]), .QN(
        my_filter_reg_coefficients_n171) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_8__11_ ( .D(
        my_filter_reg_coefficients_n425), .CK(clk), .RN(
        my_filter_reg_coefficients_n501), .Q(my_filter_q_reg_coeff[39]), .QN(
        my_filter_reg_coefficients_n172) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_8__12_ ( .D(
        my_filter_reg_coefficients_n424), .CK(clk), .RN(
        my_filter_reg_coefficients_n501), .Q(my_filter_q_reg_coeff[40]), .QN(
        my_filter_reg_coefficients_n173) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_8__13_ ( .D(
        my_filter_reg_coefficients_n423), .CK(clk), .RN(
        my_filter_reg_coefficients_n501), .Q(my_filter_q_reg_coeff[41]), .QN(
        my_filter_reg_coefficients_n174) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_7__0_ ( .D(
        my_filter_reg_coefficients_n422), .CK(clk), .RN(
        my_filter_reg_coefficients_n501), .Q(my_filter_q_reg_coeff[42]), .QN(
        my_filter_reg_coefficients_n175) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_7__1_ ( .D(
        my_filter_reg_coefficients_n421), .CK(clk), .RN(
        my_filter_reg_coefficients_n501), .Q(my_filter_q_reg_coeff[43]), .QN(
        my_filter_reg_coefficients_n176) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_7__2_ ( .D(
        my_filter_reg_coefficients_n420), .CK(clk), .RN(
        my_filter_reg_coefficients_n501), .Q(my_filter_q_reg_coeff[44]), .QN(
        my_filter_reg_coefficients_n177) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_7__3_ ( .D(
        my_filter_reg_coefficients_n419), .CK(clk), .RN(
        my_filter_reg_coefficients_n501), .Q(my_filter_q_reg_coeff[45]), .QN(
        my_filter_reg_coefficients_n178) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_7__4_ ( .D(
        my_filter_reg_coefficients_n418), .CK(clk), .RN(
        my_filter_reg_coefficients_n501), .Q(my_filter_q_reg_coeff[46]), .QN(
        my_filter_reg_coefficients_n179) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_7__5_ ( .D(
        my_filter_reg_coefficients_n417), .CK(clk), .RN(
        my_filter_reg_coefficients_n501), .Q(my_filter_q_reg_coeff[47]), .QN(
        my_filter_reg_coefficients_n180) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_7__6_ ( .D(
        my_filter_reg_coefficients_n416), .CK(clk), .RN(
        my_filter_reg_coefficients_n500), .Q(my_filter_q_reg_coeff[48]), .QN(
        my_filter_reg_coefficients_n181) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_7__7_ ( .D(
        my_filter_reg_coefficients_n415), .CK(clk), .RN(
        my_filter_reg_coefficients_n500), .Q(my_filter_q_reg_coeff[49]), .QN(
        my_filter_reg_coefficients_n182) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_7__8_ ( .D(
        my_filter_reg_coefficients_n414), .CK(clk), .RN(
        my_filter_reg_coefficients_n500), .Q(my_filter_q_reg_coeff[50]), .QN(
        my_filter_reg_coefficients_n183) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_7__9_ ( .D(
        my_filter_reg_coefficients_n413), .CK(clk), .RN(
        my_filter_reg_coefficients_n500), .Q(my_filter_q_reg_coeff[51]), .QN(
        my_filter_reg_coefficients_n184) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_7__10_ ( .D(
        my_filter_reg_coefficients_n412), .CK(clk), .RN(
        my_filter_reg_coefficients_n500), .Q(my_filter_q_reg_coeff[52]), .QN(
        my_filter_reg_coefficients_n185) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_7__11_ ( .D(
        my_filter_reg_coefficients_n411), .CK(clk), .RN(
        my_filter_reg_coefficients_n500), .Q(my_filter_q_reg_coeff[53]), .QN(
        my_filter_reg_coefficients_n186) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_7__12_ ( .D(
        my_filter_reg_coefficients_n410), .CK(clk), .RN(
        my_filter_reg_coefficients_n501), .Q(my_filter_q_reg_coeff[54]), .QN(
        my_filter_reg_coefficients_n187) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_7__13_ ( .D(
        my_filter_reg_coefficients_n409), .CK(clk), .RN(
        my_filter_reg_coefficients_n501), .Q(my_filter_q_reg_coeff[55]), .QN(
        my_filter_reg_coefficients_n188) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_6__0_ ( .D(
        my_filter_reg_coefficients_n408), .CK(clk), .RN(
        my_filter_reg_coefficients_n500), .Q(my_filter_q_reg_coeff[56]), .QN(
        my_filter_reg_coefficients_n189) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_6__1_ ( .D(
        my_filter_reg_coefficients_n407), .CK(clk), .RN(
        my_filter_reg_coefficients_n500), .Q(my_filter_q_reg_coeff[57]), .QN(
        my_filter_reg_coefficients_n190) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_6__2_ ( .D(
        my_filter_reg_coefficients_n406), .CK(clk), .RN(
        my_filter_reg_coefficients_n500), .Q(my_filter_q_reg_coeff[58]), .QN(
        my_filter_reg_coefficients_n191) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_6__3_ ( .D(
        my_filter_reg_coefficients_n405), .CK(clk), .RN(
        my_filter_reg_coefficients_n500), .Q(my_filter_q_reg_coeff[59]), .QN(
        my_filter_reg_coefficients_n192) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_6__4_ ( .D(
        my_filter_reg_coefficients_n404), .CK(clk), .RN(
        my_filter_reg_coefficients_n499), .Q(my_filter_q_reg_coeff[60]), .QN(
        my_filter_reg_coefficients_n193) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_6__5_ ( .D(
        my_filter_reg_coefficients_n403), .CK(clk), .RN(
        my_filter_reg_coefficients_n499), .Q(my_filter_q_reg_coeff[61]), .QN(
        my_filter_reg_coefficients_n194) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_6__6_ ( .D(
        my_filter_reg_coefficients_n402), .CK(clk), .RN(
        my_filter_reg_coefficients_n499), .Q(my_filter_q_reg_coeff[62]), .QN(
        my_filter_reg_coefficients_n195) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_6__7_ ( .D(
        my_filter_reg_coefficients_n401), .CK(clk), .RN(
        my_filter_reg_coefficients_n499), .Q(my_filter_q_reg_coeff[63]), .QN(
        my_filter_reg_coefficients_n196) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_6__8_ ( .D(
        my_filter_reg_coefficients_n400), .CK(clk), .RN(
        my_filter_reg_coefficients_n500), .Q(my_filter_q_reg_coeff[64]), .QN(
        my_filter_reg_coefficients_n197) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_6__9_ ( .D(
        my_filter_reg_coefficients_n399), .CK(clk), .RN(
        my_filter_reg_coefficients_n500), .Q(my_filter_q_reg_coeff[65]), .QN(
        my_filter_reg_coefficients_n198) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_6__10_ ( .D(
        my_filter_reg_coefficients_n398), .CK(clk), .RN(
        my_filter_reg_coefficients_n500), .Q(my_filter_q_reg_coeff[66]), .QN(
        my_filter_reg_coefficients_n199) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_6__11_ ( .D(
        my_filter_reg_coefficients_n397), .CK(clk), .RN(
        my_filter_reg_coefficients_n500), .Q(my_filter_q_reg_coeff[67]), .QN(
        my_filter_reg_coefficients_n200) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_6__12_ ( .D(
        my_filter_reg_coefficients_n396), .CK(clk), .RN(
        my_filter_reg_coefficients_n500), .Q(my_filter_q_reg_coeff[68]), .QN(
        my_filter_reg_coefficients_n201) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_6__13_ ( .D(
        my_filter_reg_coefficients_n395), .CK(clk), .RN(
        my_filter_reg_coefficients_n500), .Q(my_filter_q_reg_coeff[69]), .QN(
        my_filter_reg_coefficients_n202) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_5__0_ ( .D(
        my_filter_reg_coefficients_n394), .CK(clk), .RN(
        my_filter_reg_coefficients_n500), .Q(my_filter_q_reg_coeff[70]), .QN(
        my_filter_reg_coefficients_n203) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_5__1_ ( .D(
        my_filter_reg_coefficients_n393), .CK(clk), .RN(
        my_filter_reg_coefficients_n500), .Q(my_filter_q_reg_coeff[71]), .QN(
        my_filter_reg_coefficients_n204) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_5__2_ ( .D(
        my_filter_reg_coefficients_n392), .CK(clk), .RN(
        my_filter_reg_coefficients_n499), .Q(my_filter_q_reg_coeff[72]), .QN(
        my_filter_reg_coefficients_n205) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_5__3_ ( .D(
        my_filter_reg_coefficients_n391), .CK(clk), .RN(
        my_filter_reg_coefficients_n499), .Q(my_filter_q_reg_coeff[73]), .QN(
        my_filter_reg_coefficients_n206) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_5__4_ ( .D(
        my_filter_reg_coefficients_n390), .CK(clk), .RN(
        my_filter_reg_coefficients_n499), .Q(my_filter_q_reg_coeff[74]), .QN(
        my_filter_reg_coefficients_n207) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_5__5_ ( .D(
        my_filter_reg_coefficients_n389), .CK(clk), .RN(
        my_filter_reg_coefficients_n499), .Q(my_filter_q_reg_coeff[75]), .QN(
        my_filter_reg_coefficients_n208) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_5__6_ ( .D(
        my_filter_reg_coefficients_n388), .CK(clk), .RN(
        my_filter_reg_coefficients_n499), .Q(my_filter_q_reg_coeff[76]), .QN(
        my_filter_reg_coefficients_n209) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_5__7_ ( .D(
        my_filter_reg_coefficients_n387), .CK(clk), .RN(
        my_filter_reg_coefficients_n499), .Q(my_filter_q_reg_coeff[77]), .QN(
        my_filter_reg_coefficients_n210) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_5__8_ ( .D(
        my_filter_reg_coefficients_n386), .CK(clk), .RN(
        my_filter_reg_coefficients_n499), .Q(my_filter_q_reg_coeff[78]), .QN(
        my_filter_reg_coefficients_n211) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_5__9_ ( .D(
        my_filter_reg_coefficients_n385), .CK(clk), .RN(
        my_filter_reg_coefficients_n499), .Q(my_filter_q_reg_coeff[79]), .QN(
        my_filter_reg_coefficients_n212) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_5__10_ ( .D(
        my_filter_reg_coefficients_n384), .CK(clk), .RN(
        my_filter_reg_coefficients_n499), .Q(my_filter_q_reg_coeff[80]), .QN(
        my_filter_reg_coefficients_n213) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_5__11_ ( .D(
        my_filter_reg_coefficients_n383), .CK(clk), .RN(
        my_filter_reg_coefficients_n499), .Q(my_filter_q_reg_coeff[81]), .QN(
        my_filter_reg_coefficients_n214) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_5__12_ ( .D(
        my_filter_reg_coefficients_n382), .CK(clk), .RN(
        my_filter_reg_coefficients_n499), .Q(my_filter_q_reg_coeff[82]), .QN(
        my_filter_reg_coefficients_n215) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_5__13_ ( .D(
        my_filter_reg_coefficients_n381), .CK(clk), .RN(
        my_filter_reg_coefficients_n499), .Q(my_filter_q_reg_coeff[83]), .QN(
        my_filter_reg_coefficients_n216) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_4__0_ ( .D(
        my_filter_reg_coefficients_n380), .CK(clk), .RN(
        my_filter_reg_coefficients_n498), .Q(my_filter_q_reg_coeff[84]), .QN(
        my_filter_reg_coefficients_n217) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_4__1_ ( .D(
        my_filter_reg_coefficients_n379), .CK(clk), .RN(
        my_filter_reg_coefficients_n498), .Q(my_filter_q_reg_coeff[85]), .QN(
        my_filter_reg_coefficients_n218) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_4__2_ ( .D(
        my_filter_reg_coefficients_n378), .CK(clk), .RN(
        my_filter_reg_coefficients_n498), .Q(my_filter_q_reg_coeff[86]), .QN(
        my_filter_reg_coefficients_n219) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_4__3_ ( .D(
        my_filter_reg_coefficients_n377), .CK(clk), .RN(
        my_filter_reg_coefficients_n498), .Q(my_filter_q_reg_coeff[87]), .QN(
        my_filter_reg_coefficients_n220) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_4__4_ ( .D(
        my_filter_reg_coefficients_n376), .CK(clk), .RN(
        my_filter_reg_coefficients_n498), .Q(my_filter_q_reg_coeff[88]), .QN(
        my_filter_reg_coefficients_n221) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_4__5_ ( .D(
        my_filter_reg_coefficients_n375), .CK(clk), .RN(
        my_filter_reg_coefficients_n498), .Q(my_filter_q_reg_coeff[89]), .QN(
        my_filter_reg_coefficients_n222) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_4__6_ ( .D(
        my_filter_reg_coefficients_n374), .CK(clk), .RN(
        my_filter_reg_coefficients_n498), .Q(my_filter_q_reg_coeff[90]), .QN(
        my_filter_reg_coefficients_n223) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_4__7_ ( .D(
        my_filter_reg_coefficients_n373), .CK(clk), .RN(
        my_filter_reg_coefficients_n498), .Q(my_filter_q_reg_coeff[91]), .QN(
        my_filter_reg_coefficients_n224) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_4__8_ ( .D(
        my_filter_reg_coefficients_n372), .CK(clk), .RN(
        my_filter_reg_coefficients_n498), .Q(my_filter_q_reg_coeff[92]), .QN(
        my_filter_reg_coefficients_n225) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_4__9_ ( .D(
        my_filter_reg_coefficients_n371), .CK(clk), .RN(
        my_filter_reg_coefficients_n498), .Q(my_filter_q_reg_coeff[93]), .QN(
        my_filter_reg_coefficients_n226) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_4__10_ ( .D(
        my_filter_reg_coefficients_n370), .CK(clk), .RN(
        my_filter_reg_coefficients_n499), .Q(my_filter_q_reg_coeff[94]), .QN(
        my_filter_reg_coefficients_n227) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_4__11_ ( .D(
        my_filter_reg_coefficients_n369), .CK(clk), .RN(
        my_filter_reg_coefficients_n499), .Q(my_filter_q_reg_coeff[95]), .QN(
        my_filter_reg_coefficients_n228) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_4__12_ ( .D(
        my_filter_reg_coefficients_n368), .CK(clk), .RN(
        my_filter_reg_coefficients_n497), .Q(my_filter_q_reg_coeff[96]), .QN(
        my_filter_reg_coefficients_n229) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_4__13_ ( .D(
        my_filter_reg_coefficients_n367), .CK(clk), .RN(
        my_filter_reg_coefficients_n497), .Q(my_filter_q_reg_coeff[97]), .QN(
        my_filter_reg_coefficients_n230) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_3__0_ ( .D(
        my_filter_reg_coefficients_n366), .CK(clk), .RN(
        my_filter_reg_coefficients_n497), .Q(my_filter_q_reg_coeff[98]), .QN(
        my_filter_reg_coefficients_n231) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_3__1_ ( .D(
        my_filter_reg_coefficients_n365), .CK(clk), .RN(
        my_filter_reg_coefficients_n497), .Q(my_filter_q_reg_coeff[99]), .QN(
        my_filter_reg_coefficients_n232) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_3__2_ ( .D(
        my_filter_reg_coefficients_n364), .CK(clk), .RN(
        my_filter_reg_coefficients_n498), .Q(my_filter_q_reg_coeff[100]), .QN(
        my_filter_reg_coefficients_n233) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_3__3_ ( .D(
        my_filter_reg_coefficients_n363), .CK(clk), .RN(
        my_filter_reg_coefficients_n498), .Q(my_filter_q_reg_coeff[101]), .QN(
        my_filter_reg_coefficients_n234) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_3__4_ ( .D(
        my_filter_reg_coefficients_n362), .CK(clk), .RN(
        my_filter_reg_coefficients_n498), .Q(my_filter_q_reg_coeff[102]), .QN(
        my_filter_reg_coefficients_n235) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_3__5_ ( .D(
        my_filter_reg_coefficients_n361), .CK(clk), .RN(
        my_filter_reg_coefficients_n498), .Q(my_filter_q_reg_coeff[103]), .QN(
        my_filter_reg_coefficients_n236) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_3__6_ ( .D(
        my_filter_reg_coefficients_n360), .CK(clk), .RN(
        my_filter_reg_coefficients_n498), .Q(my_filter_q_reg_coeff[104]), .QN(
        my_filter_reg_coefficients_n237) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_3__7_ ( .D(
        my_filter_reg_coefficients_n359), .CK(clk), .RN(
        my_filter_reg_coefficients_n498), .Q(my_filter_q_reg_coeff[105]), .QN(
        my_filter_reg_coefficients_n238) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_3__8_ ( .D(
        my_filter_reg_coefficients_n358), .CK(clk), .RN(
        my_filter_reg_coefficients_n498), .Q(my_filter_q_reg_coeff[106]), .QN(
        my_filter_reg_coefficients_n239) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_3__9_ ( .D(
        my_filter_reg_coefficients_n357), .CK(clk), .RN(
        my_filter_reg_coefficients_n498), .Q(my_filter_q_reg_coeff[107]), .QN(
        my_filter_reg_coefficients_n240) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_3__10_ ( .D(
        my_filter_reg_coefficients_n356), .CK(clk), .RN(
        my_filter_reg_coefficients_n497), .Q(my_filter_q_reg_coeff[108]), .QN(
        my_filter_reg_coefficients_n241) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_3__11_ ( .D(
        my_filter_reg_coefficients_n355), .CK(clk), .RN(
        my_filter_reg_coefficients_n497), .Q(my_filter_q_reg_coeff[109]), .QN(
        my_filter_reg_coefficients_n242) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_3__12_ ( .D(
        my_filter_reg_coefficients_n354), .CK(clk), .RN(
        my_filter_reg_coefficients_n497), .Q(my_filter_q_reg_coeff[110]), .QN(
        my_filter_reg_coefficients_n243) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_3__13_ ( .D(
        my_filter_reg_coefficients_n353), .CK(clk), .RN(
        my_filter_reg_coefficients_n497), .Q(my_filter_q_reg_coeff[111]), .QN(
        my_filter_reg_coefficients_n244) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_2__0_ ( .D(
        my_filter_reg_coefficients_n352), .CK(clk), .RN(
        my_filter_reg_coefficients_n497), .Q(my_filter_q_reg_coeff[112]), .QN(
        my_filter_reg_coefficients_n245) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_2__1_ ( .D(
        my_filter_reg_coefficients_n351), .CK(clk), .RN(
        my_filter_reg_coefficients_n497), .Q(my_filter_q_reg_coeff[113]), .QN(
        my_filter_reg_coefficients_n246) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_2__2_ ( .D(
        my_filter_reg_coefficients_n350), .CK(clk), .RN(
        my_filter_reg_coefficients_n497), .Q(my_filter_q_reg_coeff[114]), .QN(
        my_filter_reg_coefficients_n247) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_2__3_ ( .D(
        my_filter_reg_coefficients_n349), .CK(clk), .RN(
        my_filter_reg_coefficients_n497), .Q(my_filter_q_reg_coeff[115]), .QN(
        my_filter_reg_coefficients_n248) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_2__4_ ( .D(
        my_filter_reg_coefficients_n348), .CK(clk), .RN(
        my_filter_reg_coefficients_n497), .Q(my_filter_q_reg_coeff[116]), .QN(
        my_filter_reg_coefficients_n249) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_2__5_ ( .D(
        my_filter_reg_coefficients_n347), .CK(clk), .RN(
        my_filter_reg_coefficients_n497), .Q(my_filter_q_reg_coeff[117]), .QN(
        my_filter_reg_coefficients_n250) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_2__6_ ( .D(
        my_filter_reg_coefficients_n346), .CK(clk), .RN(
        my_filter_reg_coefficients_n497), .Q(my_filter_q_reg_coeff[118]), .QN(
        my_filter_reg_coefficients_n251) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_2__7_ ( .D(
        my_filter_reg_coefficients_n345), .CK(clk), .RN(
        my_filter_reg_coefficients_n497), .Q(my_filter_q_reg_coeff[119]), .QN(
        my_filter_reg_coefficients_n252) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_2__8_ ( .D(
        my_filter_reg_coefficients_n344), .CK(clk), .RN(
        my_filter_reg_coefficients_n504), .Q(my_filter_q_reg_coeff[120]), .QN(
        my_filter_reg_coefficients_n253) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_2__9_ ( .D(
        my_filter_reg_coefficients_n343), .CK(clk), .RN(
        my_filter_reg_coefficients_n504), .Q(my_filter_q_reg_coeff[121]), .QN(
        my_filter_reg_coefficients_n254) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_2__10_ ( .D(
        my_filter_reg_coefficients_n342), .CK(clk), .RN(
        my_filter_reg_coefficients_n504), .Q(my_filter_q_reg_coeff[122]), .QN(
        my_filter_reg_coefficients_n255) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_2__11_ ( .D(
        my_filter_reg_coefficients_n341), .CK(clk), .RN(
        my_filter_reg_coefficients_n504), .Q(my_filter_q_reg_coeff[123]), .QN(
        my_filter_reg_coefficients_n256) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_2__12_ ( .D(
        my_filter_reg_coefficients_n340), .CK(clk), .RN(
        my_filter_reg_coefficients_n504), .Q(my_filter_q_reg_coeff[124]), .QN(
        my_filter_reg_coefficients_n257) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_2__13_ ( .D(
        my_filter_reg_coefficients_n339), .CK(clk), .RN(
        my_filter_reg_coefficients_n504), .Q(my_filter_q_reg_coeff[125]), .QN(
        my_filter_reg_coefficients_n258) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_1__0_ ( .D(
        my_filter_reg_coefficients_n338), .CK(clk), .RN(
        my_filter_reg_coefficients_n504), .Q(my_filter_q_reg_coeff[126]), .QN(
        my_filter_reg_coefficients_n259) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_1__1_ ( .D(
        my_filter_reg_coefficients_n337), .CK(clk), .RN(
        my_filter_reg_coefficients_n504), .Q(my_filter_q_reg_coeff[127]), .QN(
        my_filter_reg_coefficients_n260) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_1__2_ ( .D(
        my_filter_reg_coefficients_n336), .CK(clk), .RN(
        my_filter_reg_coefficients_n503), .Q(my_filter_q_reg_coeff[128]), .QN(
        my_filter_reg_coefficients_n261) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_1__3_ ( .D(
        my_filter_reg_coefficients_n335), .CK(clk), .RN(
        my_filter_reg_coefficients_n503), .Q(my_filter_q_reg_coeff[129]), .QN(
        my_filter_reg_coefficients_n262) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_1__4_ ( .D(
        my_filter_reg_coefficients_n334), .CK(clk), .RN(
        my_filter_reg_coefficients_n503), .Q(my_filter_q_reg_coeff[130]), .QN(
        my_filter_reg_coefficients_n263) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_1__5_ ( .D(
        my_filter_reg_coefficients_n333), .CK(clk), .RN(
        my_filter_reg_coefficients_n503), .Q(my_filter_q_reg_coeff[131]), .QN(
        my_filter_reg_coefficients_n264) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_1__6_ ( .D(
        my_filter_reg_coefficients_n332), .CK(clk), .RN(
        my_filter_reg_coefficients_n505), .Q(my_filter_q_reg_coeff[132]), .QN(
        my_filter_reg_coefficients_n265) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_1__7_ ( .D(
        my_filter_reg_coefficients_n331), .CK(clk), .RN(
        my_filter_reg_coefficients_n505), .Q(my_filter_q_reg_coeff[133]), .QN(
        my_filter_reg_coefficients_n266) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_1__8_ ( .D(
        my_filter_reg_coefficients_n330), .CK(clk), .RN(
        my_filter_reg_coefficients_n504), .Q(my_filter_q_reg_coeff[134]), .QN(
        my_filter_reg_coefficients_n267) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_1__9_ ( .D(
        my_filter_reg_coefficients_n329), .CK(clk), .RN(
        my_filter_reg_coefficients_n504), .Q(my_filter_q_reg_coeff[135]), .QN(
        my_filter_reg_coefficients_n268) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_1__10_ ( .D(
        my_filter_reg_coefficients_n328), .CK(clk), .RN(
        my_filter_reg_coefficients_n504), .Q(my_filter_q_reg_coeff[136]), .QN(
        my_filter_reg_coefficients_n269) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_1__11_ ( .D(
        my_filter_reg_coefficients_n327), .CK(clk), .RN(
        my_filter_reg_coefficients_n504), .Q(my_filter_q_reg_coeff[137]), .QN(
        my_filter_reg_coefficients_n270) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_1__12_ ( .D(
        my_filter_reg_coefficients_n326), .CK(clk), .RN(
        my_filter_reg_coefficients_n504), .Q(my_filter_q_reg_coeff[138]), .QN(
        my_filter_reg_coefficients_n271) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_1__13_ ( .D(
        my_filter_reg_coefficients_n325), .CK(clk), .RN(
        my_filter_reg_coefficients_n504), .Q(my_filter_q_reg_coeff[139]), .QN(
        my_filter_reg_coefficients_n272) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_0__0_ ( .D(
        my_filter_reg_coefficients_n324), .CK(clk), .RN(
        my_filter_reg_coefficients_n504), .Q(my_filter_q_reg_coeff[140]), .QN(
        my_filter_reg_coefficients_n273) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_0__1_ ( .D(
        my_filter_reg_coefficients_n323), .CK(clk), .RN(
        my_filter_reg_coefficients_n504), .Q(my_filter_q_reg_coeff[141]), .QN(
        my_filter_reg_coefficients_n274) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_0__2_ ( .D(
        my_filter_reg_coefficients_n322), .CK(clk), .RN(
        my_filter_reg_coefficients_n504), .Q(my_filter_q_reg_coeff[142]), .QN(
        my_filter_reg_coefficients_n275) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_0__3_ ( .D(
        my_filter_reg_coefficients_n321), .CK(clk), .RN(
        my_filter_reg_coefficients_n504), .Q(my_filter_q_reg_coeff[143]), .QN(
        my_filter_reg_coefficients_n276) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_0__4_ ( .D(
        my_filter_reg_coefficients_n320), .CK(clk), .RN(
        my_filter_reg_coefficients_n505), .Q(my_filter_q_reg_coeff[144]), .QN(
        my_filter_reg_coefficients_n277) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_0__5_ ( .D(
        my_filter_reg_coefficients_n319), .CK(clk), .RN(
        my_filter_reg_coefficients_n505), .Q(my_filter_q_reg_coeff[145]), .QN(
        my_filter_reg_coefficients_n278) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_0__6_ ( .D(
        my_filter_reg_coefficients_n318), .CK(clk), .RN(
        my_filter_reg_coefficients_n505), .Q(my_filter_q_reg_coeff[146]), .QN(
        my_filter_reg_coefficients_n279) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_0__7_ ( .D(
        my_filter_reg_coefficients_n317), .CK(clk), .RN(
        my_filter_reg_coefficients_n505), .Q(my_filter_q_reg_coeff[147]), .QN(
        my_filter_reg_coefficients_n280) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_0__8_ ( .D(
        my_filter_reg_coefficients_n316), .CK(clk), .RN(
        my_filter_reg_coefficients_n505), .Q(my_filter_q_reg_coeff[148]), .QN(
        my_filter_reg_coefficients_n281) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_0__9_ ( .D(
        my_filter_reg_coefficients_n315), .CK(clk), .RN(
        my_filter_reg_coefficients_n505), .Q(my_filter_q_reg_coeff[149]), .QN(
        my_filter_reg_coefficients_n282) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_0__10_ ( .D(
        my_filter_reg_coefficients_n314), .CK(clk), .RN(
        my_filter_reg_coefficients_n505), .Q(my_filter_q_reg_coeff[150]), .QN(
        my_filter_reg_coefficients_n283) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_0__11_ ( .D(
        my_filter_reg_coefficients_n313), .CK(clk), .RN(
        my_filter_reg_coefficients_n505), .Q(my_filter_q_reg_coeff[151]), .QN(
        my_filter_reg_coefficients_n284) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_0__12_ ( .D(
        my_filter_reg_coefficients_n312), .CK(clk), .RN(
        my_filter_reg_coefficients_n505), .Q(my_filter_q_reg_coeff[152]), .QN(
        my_filter_reg_coefficients_n285) );
  DFFR_X1 my_filter_reg_coefficients_q_reg_0__13_ ( .D(
        my_filter_reg_coefficients_n311), .CK(clk), .RN(
        my_filter_reg_coefficients_n505), .Q(my_filter_q_reg_coeff[153]), .QN(
        my_filter_reg_coefficients_n286) );
  INV_X1 my_filter_reg_out_U33 ( .A(my_filter_en_reg_out), .ZN(
        my_filter_reg_out_n47) );
  NAND2_X1 my_filter_reg_out_U32 ( .A1(my_filter_reg_out_n46), .A2(
        my_filter_reg_out_n47), .ZN(my_filter_reg_out_n2) );
  NAND2_X1 my_filter_reg_out_U31 ( .A1(my_filter_data_sum[0]), .A2(
        my_filter_en_reg_out), .ZN(my_filter_reg_out_n16) );
  OAI21_X1 my_filter_reg_out_U30 ( .B1(my_filter_reg_out_n2), .B2(
        my_filter_reg_out_n27), .A(my_filter_reg_out_n16), .ZN(
        my_filter_reg_out_n44) );
  NAND2_X1 my_filter_reg_out_U29 ( .A1(my_filter_data_sum[5]), .A2(
        my_filter_en_reg_out), .ZN(my_filter_reg_out_n11) );
  OAI21_X1 my_filter_reg_out_U28 ( .B1(my_filter_reg_out_n2), .B2(
        my_filter_reg_out_n17), .A(my_filter_reg_out_n11), .ZN(
        my_filter_reg_out_n39) );
  NAND2_X1 my_filter_reg_out_U27 ( .A1(my_filter_data_sum[4]), .A2(
        my_filter_en_reg_out), .ZN(my_filter_reg_out_n12) );
  OAI21_X1 my_filter_reg_out_U26 ( .B1(my_filter_reg_out_n2), .B2(
        my_filter_reg_out_n30), .A(my_filter_reg_out_n12), .ZN(
        my_filter_reg_out_n40) );
  NAND2_X1 my_filter_reg_out_U25 ( .A1(my_filter_data_sum[3]), .A2(
        my_filter_en_reg_out), .ZN(my_filter_reg_out_n13) );
  OAI21_X1 my_filter_reg_out_U24 ( .B1(my_filter_reg_out_n2), .B2(
        my_filter_reg_out_n29), .A(my_filter_reg_out_n13), .ZN(
        my_filter_reg_out_n41) );
  NAND2_X1 my_filter_reg_out_U23 ( .A1(my_filter_data_sum[2]), .A2(
        my_filter_en_reg_out), .ZN(my_filter_reg_out_n14) );
  OAI21_X1 my_filter_reg_out_U22 ( .B1(my_filter_reg_out_n2), .B2(
        my_filter_reg_out_n28), .A(my_filter_reg_out_n14), .ZN(
        my_filter_reg_out_n42) );
  NAND2_X1 my_filter_reg_out_U21 ( .A1(my_filter_data_sum[1]), .A2(
        my_filter_en_reg_out), .ZN(my_filter_reg_out_n15) );
  OAI21_X1 my_filter_reg_out_U20 ( .B1(my_filter_reg_out_n2), .B2(
        my_filter_reg_out_n26), .A(my_filter_reg_out_n15), .ZN(
        my_filter_reg_out_n43) );
  NAND2_X1 my_filter_reg_out_U19 ( .A1(my_filter_en_reg_out), .A2(
        my_filter_data_sum[13]), .ZN(my_filter_reg_out_n3) );
  OAI21_X1 my_filter_reg_out_U18 ( .B1(my_filter_reg_out_n2), .B2(
        my_filter_reg_out_n25), .A(my_filter_reg_out_n3), .ZN(
        my_filter_reg_out_n31) );
  NAND2_X1 my_filter_reg_out_U17 ( .A1(my_filter_data_sum[12]), .A2(
        my_filter_en_reg_out), .ZN(my_filter_reg_out_n4) );
  OAI21_X1 my_filter_reg_out_U16 ( .B1(my_filter_reg_out_n2), .B2(
        my_filter_reg_out_n24), .A(my_filter_reg_out_n4), .ZN(
        my_filter_reg_out_n32) );
  NAND2_X1 my_filter_reg_out_U15 ( .A1(my_filter_data_sum[11]), .A2(
        my_filter_en_reg_out), .ZN(my_filter_reg_out_n5) );
  OAI21_X1 my_filter_reg_out_U14 ( .B1(my_filter_reg_out_n2), .B2(
        my_filter_reg_out_n23), .A(my_filter_reg_out_n5), .ZN(
        my_filter_reg_out_n33) );
  NAND2_X1 my_filter_reg_out_U13 ( .A1(my_filter_data_sum[10]), .A2(
        my_filter_en_reg_out), .ZN(my_filter_reg_out_n6) );
  OAI21_X1 my_filter_reg_out_U12 ( .B1(my_filter_reg_out_n2), .B2(
        my_filter_reg_out_n22), .A(my_filter_reg_out_n6), .ZN(
        my_filter_reg_out_n34) );
  NAND2_X1 my_filter_reg_out_U11 ( .A1(my_filter_data_sum[9]), .A2(
        my_filter_en_reg_out), .ZN(my_filter_reg_out_n7) );
  OAI21_X1 my_filter_reg_out_U10 ( .B1(my_filter_reg_out_n2), .B2(
        my_filter_reg_out_n21), .A(my_filter_reg_out_n7), .ZN(
        my_filter_reg_out_n35) );
  NAND2_X1 my_filter_reg_out_U9 ( .A1(my_filter_data_sum[8]), .A2(
        my_filter_en_reg_out), .ZN(my_filter_reg_out_n8) );
  OAI21_X1 my_filter_reg_out_U8 ( .B1(my_filter_reg_out_n2), .B2(
        my_filter_reg_out_n20), .A(my_filter_reg_out_n8), .ZN(
        my_filter_reg_out_n36) );
  NAND2_X1 my_filter_reg_out_U7 ( .A1(my_filter_data_sum[7]), .A2(
        my_filter_en_reg_out), .ZN(my_filter_reg_out_n9) );
  OAI21_X1 my_filter_reg_out_U6 ( .B1(my_filter_reg_out_n2), .B2(
        my_filter_reg_out_n19), .A(my_filter_reg_out_n9), .ZN(
        my_filter_reg_out_n37) );
  NAND2_X1 my_filter_reg_out_U5 ( .A1(my_filter_data_sum[6]), .A2(
        my_filter_en_reg_out), .ZN(my_filter_reg_out_n10) );
  OAI21_X1 my_filter_reg_out_U4 ( .B1(my_filter_reg_out_n2), .B2(
        my_filter_reg_out_n18), .A(my_filter_reg_out_n10), .ZN(
        my_filter_reg_out_n38) );
  BUF_X1 my_filter_reg_out_U3 ( .A(my_filter_n2), .Z(my_filter_reg_out_n46) );
  DFFR_X1 my_filter_reg_out_q_reg_0_ ( .D(my_filter_reg_out_n44), .CK(clk), 
        .RN(my_filter_reg_out_n46), .Q(dout[0]), .QN(my_filter_reg_out_n27) );
  DFFR_X1 my_filter_reg_out_q_reg_1_ ( .D(my_filter_reg_out_n43), .CK(clk), 
        .RN(my_filter_reg_out_n46), .Q(dout[1]), .QN(my_filter_reg_out_n26) );
  DFFR_X1 my_filter_reg_out_q_reg_2_ ( .D(my_filter_reg_out_n42), .CK(clk), 
        .RN(my_filter_reg_out_n46), .Q(dout[2]), .QN(my_filter_reg_out_n28) );
  DFFR_X1 my_filter_reg_out_q_reg_3_ ( .D(my_filter_reg_out_n41), .CK(clk), 
        .RN(my_filter_reg_out_n46), .Q(dout[3]), .QN(my_filter_reg_out_n29) );
  DFFR_X1 my_filter_reg_out_q_reg_4_ ( .D(my_filter_reg_out_n40), .CK(clk), 
        .RN(my_filter_reg_out_n46), .Q(dout[4]), .QN(my_filter_reg_out_n30) );
  DFFR_X1 my_filter_reg_out_q_reg_5_ ( .D(my_filter_reg_out_n39), .CK(clk), 
        .RN(my_filter_reg_out_n46), .Q(dout[5]), .QN(my_filter_reg_out_n17) );
  DFFR_X1 my_filter_reg_out_q_reg_6_ ( .D(my_filter_reg_out_n38), .CK(clk), 
        .RN(my_filter_reg_out_n46), .Q(dout[6]), .QN(my_filter_reg_out_n18) );
  DFFR_X1 my_filter_reg_out_q_reg_7_ ( .D(my_filter_reg_out_n37), .CK(clk), 
        .RN(my_filter_reg_out_n46), .Q(dout[7]), .QN(my_filter_reg_out_n19) );
  DFFR_X1 my_filter_reg_out_q_reg_8_ ( .D(my_filter_reg_out_n36), .CK(clk), 
        .RN(my_filter_reg_out_n46), .Q(dout[8]), .QN(my_filter_reg_out_n20) );
  DFFR_X1 my_filter_reg_out_q_reg_9_ ( .D(my_filter_reg_out_n35), .CK(clk), 
        .RN(my_filter_reg_out_n46), .Q(dout[9]), .QN(my_filter_reg_out_n21) );
  DFFR_X1 my_filter_reg_out_q_reg_10_ ( .D(my_filter_reg_out_n34), .CK(clk), 
        .RN(my_filter_reg_out_n46), .Q(dout[10]), .QN(my_filter_reg_out_n22)
         );
  DFFR_X1 my_filter_reg_out_q_reg_11_ ( .D(my_filter_reg_out_n33), .CK(clk), 
        .RN(my_filter_reg_out_n46), .Q(dout[11]), .QN(my_filter_reg_out_n23)
         );
  DFFR_X1 my_filter_reg_out_q_reg_12_ ( .D(my_filter_reg_out_n32), .CK(clk), 
        .RN(my_filter_reg_out_n46), .Q(dout[12]), .QN(my_filter_reg_out_n24)
         );
  DFFR_X1 my_filter_reg_out_q_reg_13_ ( .D(my_filter_reg_out_n31), .CK(clk), 
        .RN(my_filter_reg_out_n46), .Q(dout[13]), .QN(my_filter_reg_out_n25)
         );
  DFFR_X1 my_filter_ff_en_reg_out_q_reg ( .D(vin), .CK(clk), .RN(my_filter_n2), 
        .Q(my_filter_en_reg_out) );
  DFFR_X1 my_filter_ff_vout_q_reg ( .D(my_filter_en_reg_out), .CK(clk), .RN(
        my_filter_n2), .Q(vout) );
  BUF_X1 my_filter_delay_line_U8 ( .A(vin), .Z(my_filter_delay_line_n8) );
  BUF_X1 my_filter_delay_line_U7 ( .A(my_filter_n2), .Z(
        my_filter_delay_line_n10) );
  BUF_X1 my_filter_delay_line_U6 ( .A(my_filter_n2), .Z(
        my_filter_delay_line_n9) );
  BUF_X1 my_filter_delay_line_U5 ( .A(my_filter_delay_line_n10), .Z(
        my_filter_delay_line_n15) );
  BUF_X1 my_filter_delay_line_U4 ( .A(my_filter_delay_line_n10), .Z(
        my_filter_delay_line_n14) );
  BUF_X1 my_filter_delay_line_U3 ( .A(my_filter_delay_line_n9), .Z(
        my_filter_delay_line_n13) );
  BUF_X1 my_filter_delay_line_U2 ( .A(my_filter_delay_line_n9), .Z(
        my_filter_delay_line_n12) );
  BUF_X1 my_filter_delay_line_U1 ( .A(my_filter_delay_line_n9), .Z(
        my_filter_delay_line_n11) );
  NAND2_X1 my_filter_delay_line_delay_chain_0_U34 ( .A1(
        my_filter_delay_line_n8), .A2(my_filter_q_reg_samp_13_), .ZN(
        my_filter_delay_line_delay_chain_0_n3) );
  OAI21_X1 my_filter_delay_line_delay_chain_0_U33 ( .B1(
        my_filter_delay_line_delay_chain_0_n2), .B2(
        my_filter_delay_line_delay_chain_0_n30), .A(
        my_filter_delay_line_delay_chain_0_n3), .ZN(
        my_filter_delay_line_delay_chain_0_n31) );
  NAND2_X1 my_filter_delay_line_delay_chain_0_U32 ( .A1(
        my_filter_q_reg_samp_12_), .A2(my_filter_delay_line_n8), .ZN(
        my_filter_delay_line_delay_chain_0_n4) );
  OAI21_X1 my_filter_delay_line_delay_chain_0_U31 ( .B1(
        my_filter_delay_line_delay_chain_0_n2), .B2(
        my_filter_delay_line_delay_chain_0_n29), .A(
        my_filter_delay_line_delay_chain_0_n4), .ZN(
        my_filter_delay_line_delay_chain_0_n32) );
  NAND2_X1 my_filter_delay_line_delay_chain_0_U30 ( .A1(
        my_filter_q_reg_samp_11_), .A2(my_filter_delay_line_delay_chain_0_n48), 
        .ZN(my_filter_delay_line_delay_chain_0_n5) );
  OAI21_X1 my_filter_delay_line_delay_chain_0_U29 ( .B1(
        my_filter_delay_line_delay_chain_0_n2), .B2(
        my_filter_delay_line_delay_chain_0_n28), .A(
        my_filter_delay_line_delay_chain_0_n5), .ZN(
        my_filter_delay_line_delay_chain_0_n33) );
  NAND2_X1 my_filter_delay_line_delay_chain_0_U28 ( .A1(
        my_filter_q_reg_samp_10_), .A2(my_filter_delay_line_delay_chain_0_n48), 
        .ZN(my_filter_delay_line_delay_chain_0_n6) );
  OAI21_X1 my_filter_delay_line_delay_chain_0_U27 ( .B1(
        my_filter_delay_line_delay_chain_0_n2), .B2(
        my_filter_delay_line_delay_chain_0_n27), .A(
        my_filter_delay_line_delay_chain_0_n6), .ZN(
        my_filter_delay_line_delay_chain_0_n34) );
  NAND2_X1 my_filter_delay_line_delay_chain_0_U26 ( .A1(
        my_filter_q_reg_samp_9_), .A2(my_filter_delay_line_delay_chain_0_n48), 
        .ZN(my_filter_delay_line_delay_chain_0_n7) );
  OAI21_X1 my_filter_delay_line_delay_chain_0_U25 ( .B1(
        my_filter_delay_line_delay_chain_0_n2), .B2(
        my_filter_delay_line_delay_chain_0_n26), .A(
        my_filter_delay_line_delay_chain_0_n7), .ZN(
        my_filter_delay_line_delay_chain_0_n35) );
  NAND2_X1 my_filter_delay_line_delay_chain_0_U24 ( .A1(
        my_filter_q_reg_samp_8_), .A2(my_filter_delay_line_delay_chain_0_n48), 
        .ZN(my_filter_delay_line_delay_chain_0_n8) );
  OAI21_X1 my_filter_delay_line_delay_chain_0_U23 ( .B1(
        my_filter_delay_line_delay_chain_0_n2), .B2(
        my_filter_delay_line_delay_chain_0_n25), .A(
        my_filter_delay_line_delay_chain_0_n8), .ZN(
        my_filter_delay_line_delay_chain_0_n36) );
  NAND2_X1 my_filter_delay_line_delay_chain_0_U22 ( .A1(
        my_filter_q_reg_samp_7_), .A2(my_filter_delay_line_delay_chain_0_n48), 
        .ZN(my_filter_delay_line_delay_chain_0_n9) );
  OAI21_X1 my_filter_delay_line_delay_chain_0_U21 ( .B1(
        my_filter_delay_line_delay_chain_0_n2), .B2(
        my_filter_delay_line_delay_chain_0_n24), .A(
        my_filter_delay_line_delay_chain_0_n9), .ZN(
        my_filter_delay_line_delay_chain_0_n37) );
  NAND2_X1 my_filter_delay_line_delay_chain_0_U20 ( .A1(
        my_filter_q_reg_samp_6_), .A2(my_filter_delay_line_delay_chain_0_n48), 
        .ZN(my_filter_delay_line_delay_chain_0_n10) );
  OAI21_X1 my_filter_delay_line_delay_chain_0_U19 ( .B1(
        my_filter_delay_line_delay_chain_0_n2), .B2(
        my_filter_delay_line_delay_chain_0_n23), .A(
        my_filter_delay_line_delay_chain_0_n10), .ZN(
        my_filter_delay_line_delay_chain_0_n38) );
  NAND2_X1 my_filter_delay_line_delay_chain_0_U18 ( .A1(
        my_filter_q_reg_samp_5_), .A2(my_filter_delay_line_delay_chain_0_n48), 
        .ZN(my_filter_delay_line_delay_chain_0_n11) );
  OAI21_X1 my_filter_delay_line_delay_chain_0_U17 ( .B1(
        my_filter_delay_line_delay_chain_0_n2), .B2(
        my_filter_delay_line_delay_chain_0_n22), .A(
        my_filter_delay_line_delay_chain_0_n11), .ZN(
        my_filter_delay_line_delay_chain_0_n39) );
  NAND2_X1 my_filter_delay_line_delay_chain_0_U16 ( .A1(
        my_filter_q_reg_samp_4_), .A2(my_filter_delay_line_delay_chain_0_n48), 
        .ZN(my_filter_delay_line_delay_chain_0_n12) );
  OAI21_X1 my_filter_delay_line_delay_chain_0_U15 ( .B1(
        my_filter_delay_line_delay_chain_0_n2), .B2(
        my_filter_delay_line_delay_chain_0_n21), .A(
        my_filter_delay_line_delay_chain_0_n12), .ZN(
        my_filter_delay_line_delay_chain_0_n40) );
  NAND2_X1 my_filter_delay_line_delay_chain_0_U14 ( .A1(
        my_filter_q_reg_samp_3_), .A2(my_filter_delay_line_delay_chain_0_n48), 
        .ZN(my_filter_delay_line_delay_chain_0_n13) );
  OAI21_X1 my_filter_delay_line_delay_chain_0_U13 ( .B1(
        my_filter_delay_line_delay_chain_0_n2), .B2(
        my_filter_delay_line_delay_chain_0_n20), .A(
        my_filter_delay_line_delay_chain_0_n13), .ZN(
        my_filter_delay_line_delay_chain_0_n41) );
  NAND2_X1 my_filter_delay_line_delay_chain_0_U12 ( .A1(
        my_filter_q_reg_samp_2_), .A2(my_filter_delay_line_delay_chain_0_n48), 
        .ZN(my_filter_delay_line_delay_chain_0_n14) );
  OAI21_X1 my_filter_delay_line_delay_chain_0_U11 ( .B1(
        my_filter_delay_line_delay_chain_0_n2), .B2(
        my_filter_delay_line_delay_chain_0_n19), .A(
        my_filter_delay_line_delay_chain_0_n14), .ZN(
        my_filter_delay_line_delay_chain_0_n42) );
  NAND2_X1 my_filter_delay_line_delay_chain_0_U10 ( .A1(
        my_filter_q_reg_samp_1_), .A2(my_filter_delay_line_delay_chain_0_n48), 
        .ZN(my_filter_delay_line_delay_chain_0_n15) );
  OAI21_X1 my_filter_delay_line_delay_chain_0_U9 ( .B1(
        my_filter_delay_line_delay_chain_0_n2), .B2(
        my_filter_delay_line_delay_chain_0_n18), .A(
        my_filter_delay_line_delay_chain_0_n15), .ZN(
        my_filter_delay_line_delay_chain_0_n43) );
  NAND2_X1 my_filter_delay_line_delay_chain_0_U8 ( .A1(my_filter_q_reg_samp_0_), .A2(my_filter_delay_line_delay_chain_0_n48), .ZN(
        my_filter_delay_line_delay_chain_0_n16) );
  OAI21_X1 my_filter_delay_line_delay_chain_0_U7 ( .B1(
        my_filter_delay_line_delay_chain_0_n2), .B2(
        my_filter_delay_line_delay_chain_0_n17), .A(
        my_filter_delay_line_delay_chain_0_n16), .ZN(
        my_filter_delay_line_delay_chain_0_n44) );
  INV_X1 my_filter_delay_line_delay_chain_0_U6 ( .A(my_filter_delay_line_n8), 
        .ZN(my_filter_delay_line_delay_chain_0_n49) );
  INV_X1 my_filter_delay_line_delay_chain_0_U5 ( .A(
        my_filter_delay_line_delay_chain_0_n49), .ZN(
        my_filter_delay_line_delay_chain_0_n48) );
  NAND2_X1 my_filter_delay_line_delay_chain_0_U4 ( .A1(
        my_filter_delay_line_delay_chain_0_n50), .A2(
        my_filter_delay_line_delay_chain_0_n49), .ZN(
        my_filter_delay_line_delay_chain_0_n2) );
  BUF_X1 my_filter_delay_line_delay_chain_0_U3 ( .A(my_filter_delay_line_n15), 
        .Z(my_filter_delay_line_delay_chain_0_n50) );
  DFFR_X1 my_filter_delay_line_delay_chain_0_q_reg_0_ ( .D(
        my_filter_delay_line_delay_chain_0_n44), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_0_n50), .Q(
        my_filter_q_reg_chain_1__0_), .QN(
        my_filter_delay_line_delay_chain_0_n17) );
  DFFR_X1 my_filter_delay_line_delay_chain_0_q_reg_1_ ( .D(
        my_filter_delay_line_delay_chain_0_n43), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_0_n50), .Q(
        my_filter_q_reg_chain_1__1_), .QN(
        my_filter_delay_line_delay_chain_0_n18) );
  DFFR_X1 my_filter_delay_line_delay_chain_0_q_reg_2_ ( .D(
        my_filter_delay_line_delay_chain_0_n42), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_0_n50), .Q(
        my_filter_q_reg_chain_1__2_), .QN(
        my_filter_delay_line_delay_chain_0_n19) );
  DFFR_X1 my_filter_delay_line_delay_chain_0_q_reg_3_ ( .D(
        my_filter_delay_line_delay_chain_0_n41), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_0_n50), .Q(
        my_filter_q_reg_chain_1__3_), .QN(
        my_filter_delay_line_delay_chain_0_n20) );
  DFFR_X1 my_filter_delay_line_delay_chain_0_q_reg_4_ ( .D(
        my_filter_delay_line_delay_chain_0_n40), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_0_n50), .Q(
        my_filter_q_reg_chain_1__4_), .QN(
        my_filter_delay_line_delay_chain_0_n21) );
  DFFR_X1 my_filter_delay_line_delay_chain_0_q_reg_5_ ( .D(
        my_filter_delay_line_delay_chain_0_n39), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_0_n50), .Q(
        my_filter_q_reg_chain_1__5_), .QN(
        my_filter_delay_line_delay_chain_0_n22) );
  DFFR_X1 my_filter_delay_line_delay_chain_0_q_reg_6_ ( .D(
        my_filter_delay_line_delay_chain_0_n38), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_0_n50), .Q(
        my_filter_q_reg_chain_1__6_), .QN(
        my_filter_delay_line_delay_chain_0_n23) );
  DFFR_X1 my_filter_delay_line_delay_chain_0_q_reg_7_ ( .D(
        my_filter_delay_line_delay_chain_0_n37), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_0_n50), .Q(
        my_filter_q_reg_chain_1__7_), .QN(
        my_filter_delay_line_delay_chain_0_n24) );
  DFFR_X1 my_filter_delay_line_delay_chain_0_q_reg_8_ ( .D(
        my_filter_delay_line_delay_chain_0_n36), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_0_n50), .Q(
        my_filter_q_reg_chain_1__8_), .QN(
        my_filter_delay_line_delay_chain_0_n25) );
  DFFR_X1 my_filter_delay_line_delay_chain_0_q_reg_9_ ( .D(
        my_filter_delay_line_delay_chain_0_n35), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_0_n50), .Q(
        my_filter_q_reg_chain_1__9_), .QN(
        my_filter_delay_line_delay_chain_0_n26) );
  DFFR_X1 my_filter_delay_line_delay_chain_0_q_reg_10_ ( .D(
        my_filter_delay_line_delay_chain_0_n34), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_0_n50), .Q(
        my_filter_q_reg_chain_1__10_), .QN(
        my_filter_delay_line_delay_chain_0_n27) );
  DFFR_X1 my_filter_delay_line_delay_chain_0_q_reg_11_ ( .D(
        my_filter_delay_line_delay_chain_0_n33), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_0_n50), .Q(
        my_filter_q_reg_chain_1__11_), .QN(
        my_filter_delay_line_delay_chain_0_n28) );
  DFFR_X1 my_filter_delay_line_delay_chain_0_q_reg_12_ ( .D(
        my_filter_delay_line_delay_chain_0_n32), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_0_n50), .Q(
        my_filter_q_reg_chain_1__12_), .QN(
        my_filter_delay_line_delay_chain_0_n29) );
  DFFR_X1 my_filter_delay_line_delay_chain_0_q_reg_13_ ( .D(
        my_filter_delay_line_delay_chain_0_n31), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_0_n50), .Q(
        my_filter_q_reg_chain_1__13_), .QN(
        my_filter_delay_line_delay_chain_0_n30) );
  INV_X1 my_filter_delay_line_delay_chain_1_U35 ( .A(
        my_filter_delay_line_delay_chain_1_n50), .ZN(
        my_filter_delay_line_delay_chain_1_n49) );
  NAND2_X1 my_filter_delay_line_delay_chain_1_U34 ( .A1(
        my_filter_delay_line_delay_chain_1_n49), .A2(
        my_filter_q_reg_chain_1__13_), .ZN(
        my_filter_delay_line_delay_chain_1_n93) );
  OAI21_X1 my_filter_delay_line_delay_chain_1_U33 ( .B1(
        my_filter_delay_line_delay_chain_1_n94), .B2(
        my_filter_delay_line_delay_chain_1_n66), .A(
        my_filter_delay_line_delay_chain_1_n93), .ZN(
        my_filter_delay_line_delay_chain_1_n65) );
  NAND2_X1 my_filter_delay_line_delay_chain_1_U32 ( .A1(
        my_filter_q_reg_chain_1__12_), .A2(
        my_filter_delay_line_delay_chain_1_n49), .ZN(
        my_filter_delay_line_delay_chain_1_n92) );
  OAI21_X1 my_filter_delay_line_delay_chain_1_U31 ( .B1(
        my_filter_delay_line_delay_chain_1_n94), .B2(
        my_filter_delay_line_delay_chain_1_n67), .A(
        my_filter_delay_line_delay_chain_1_n92), .ZN(
        my_filter_delay_line_delay_chain_1_n64) );
  NAND2_X1 my_filter_delay_line_delay_chain_1_U30 ( .A1(
        my_filter_q_reg_chain_1__11_), .A2(
        my_filter_delay_line_delay_chain_1_n48), .ZN(
        my_filter_delay_line_delay_chain_1_n91) );
  OAI21_X1 my_filter_delay_line_delay_chain_1_U29 ( .B1(
        my_filter_delay_line_delay_chain_1_n94), .B2(
        my_filter_delay_line_delay_chain_1_n68), .A(
        my_filter_delay_line_delay_chain_1_n91), .ZN(
        my_filter_delay_line_delay_chain_1_n63) );
  NAND2_X1 my_filter_delay_line_delay_chain_1_U28 ( .A1(
        my_filter_q_reg_chain_1__10_), .A2(
        my_filter_delay_line_delay_chain_1_n48), .ZN(
        my_filter_delay_line_delay_chain_1_n90) );
  OAI21_X1 my_filter_delay_line_delay_chain_1_U27 ( .B1(
        my_filter_delay_line_delay_chain_1_n94), .B2(
        my_filter_delay_line_delay_chain_1_n69), .A(
        my_filter_delay_line_delay_chain_1_n90), .ZN(
        my_filter_delay_line_delay_chain_1_n62) );
  NAND2_X1 my_filter_delay_line_delay_chain_1_U26 ( .A1(
        my_filter_q_reg_chain_1__9_), .A2(
        my_filter_delay_line_delay_chain_1_n48), .ZN(
        my_filter_delay_line_delay_chain_1_n89) );
  OAI21_X1 my_filter_delay_line_delay_chain_1_U25 ( .B1(
        my_filter_delay_line_delay_chain_1_n94), .B2(
        my_filter_delay_line_delay_chain_1_n70), .A(
        my_filter_delay_line_delay_chain_1_n89), .ZN(
        my_filter_delay_line_delay_chain_1_n61) );
  NAND2_X1 my_filter_delay_line_delay_chain_1_U24 ( .A1(
        my_filter_q_reg_chain_1__8_), .A2(
        my_filter_delay_line_delay_chain_1_n48), .ZN(
        my_filter_delay_line_delay_chain_1_n88) );
  OAI21_X1 my_filter_delay_line_delay_chain_1_U23 ( .B1(
        my_filter_delay_line_delay_chain_1_n94), .B2(
        my_filter_delay_line_delay_chain_1_n71), .A(
        my_filter_delay_line_delay_chain_1_n88), .ZN(
        my_filter_delay_line_delay_chain_1_n60) );
  NAND2_X1 my_filter_delay_line_delay_chain_1_U22 ( .A1(
        my_filter_q_reg_chain_1__7_), .A2(
        my_filter_delay_line_delay_chain_1_n48), .ZN(
        my_filter_delay_line_delay_chain_1_n87) );
  OAI21_X1 my_filter_delay_line_delay_chain_1_U21 ( .B1(
        my_filter_delay_line_delay_chain_1_n94), .B2(
        my_filter_delay_line_delay_chain_1_n72), .A(
        my_filter_delay_line_delay_chain_1_n87), .ZN(
        my_filter_delay_line_delay_chain_1_n59) );
  NAND2_X1 my_filter_delay_line_delay_chain_1_U20 ( .A1(
        my_filter_q_reg_chain_1__6_), .A2(
        my_filter_delay_line_delay_chain_1_n48), .ZN(
        my_filter_delay_line_delay_chain_1_n86) );
  OAI21_X1 my_filter_delay_line_delay_chain_1_U19 ( .B1(
        my_filter_delay_line_delay_chain_1_n94), .B2(
        my_filter_delay_line_delay_chain_1_n73), .A(
        my_filter_delay_line_delay_chain_1_n86), .ZN(
        my_filter_delay_line_delay_chain_1_n58) );
  NAND2_X1 my_filter_delay_line_delay_chain_1_U18 ( .A1(
        my_filter_q_reg_chain_1__5_), .A2(
        my_filter_delay_line_delay_chain_1_n48), .ZN(
        my_filter_delay_line_delay_chain_1_n85) );
  OAI21_X1 my_filter_delay_line_delay_chain_1_U17 ( .B1(
        my_filter_delay_line_delay_chain_1_n94), .B2(
        my_filter_delay_line_delay_chain_1_n74), .A(
        my_filter_delay_line_delay_chain_1_n85), .ZN(
        my_filter_delay_line_delay_chain_1_n57) );
  NAND2_X1 my_filter_delay_line_delay_chain_1_U16 ( .A1(
        my_filter_q_reg_chain_1__4_), .A2(
        my_filter_delay_line_delay_chain_1_n48), .ZN(
        my_filter_delay_line_delay_chain_1_n84) );
  OAI21_X1 my_filter_delay_line_delay_chain_1_U15 ( .B1(
        my_filter_delay_line_delay_chain_1_n94), .B2(
        my_filter_delay_line_delay_chain_1_n75), .A(
        my_filter_delay_line_delay_chain_1_n84), .ZN(
        my_filter_delay_line_delay_chain_1_n56) );
  NAND2_X1 my_filter_delay_line_delay_chain_1_U14 ( .A1(
        my_filter_q_reg_chain_1__3_), .A2(
        my_filter_delay_line_delay_chain_1_n48), .ZN(
        my_filter_delay_line_delay_chain_1_n83) );
  OAI21_X1 my_filter_delay_line_delay_chain_1_U13 ( .B1(
        my_filter_delay_line_delay_chain_1_n94), .B2(
        my_filter_delay_line_delay_chain_1_n76), .A(
        my_filter_delay_line_delay_chain_1_n83), .ZN(
        my_filter_delay_line_delay_chain_1_n55) );
  NAND2_X1 my_filter_delay_line_delay_chain_1_U12 ( .A1(
        my_filter_q_reg_chain_1__2_), .A2(
        my_filter_delay_line_delay_chain_1_n48), .ZN(
        my_filter_delay_line_delay_chain_1_n82) );
  OAI21_X1 my_filter_delay_line_delay_chain_1_U11 ( .B1(
        my_filter_delay_line_delay_chain_1_n94), .B2(
        my_filter_delay_line_delay_chain_1_n77), .A(
        my_filter_delay_line_delay_chain_1_n82), .ZN(
        my_filter_delay_line_delay_chain_1_n54) );
  NAND2_X1 my_filter_delay_line_delay_chain_1_U10 ( .A1(
        my_filter_q_reg_chain_1__1_), .A2(
        my_filter_delay_line_delay_chain_1_n48), .ZN(
        my_filter_delay_line_delay_chain_1_n81) );
  OAI21_X1 my_filter_delay_line_delay_chain_1_U9 ( .B1(
        my_filter_delay_line_delay_chain_1_n94), .B2(
        my_filter_delay_line_delay_chain_1_n78), .A(
        my_filter_delay_line_delay_chain_1_n81), .ZN(
        my_filter_delay_line_delay_chain_1_n53) );
  NAND2_X1 my_filter_delay_line_delay_chain_1_U8 ( .A1(
        my_filter_q_reg_chain_1__0_), .A2(
        my_filter_delay_line_delay_chain_1_n48), .ZN(
        my_filter_delay_line_delay_chain_1_n80) );
  OAI21_X1 my_filter_delay_line_delay_chain_1_U7 ( .B1(
        my_filter_delay_line_delay_chain_1_n94), .B2(
        my_filter_delay_line_delay_chain_1_n79), .A(
        my_filter_delay_line_delay_chain_1_n80), .ZN(
        my_filter_delay_line_delay_chain_1_n52) );
  INV_X1 my_filter_delay_line_delay_chain_1_U6 ( .A(my_filter_delay_line_n8), 
        .ZN(my_filter_delay_line_delay_chain_1_n50) );
  INV_X1 my_filter_delay_line_delay_chain_1_U5 ( .A(
        my_filter_delay_line_delay_chain_1_n50), .ZN(
        my_filter_delay_line_delay_chain_1_n48) );
  NAND2_X1 my_filter_delay_line_delay_chain_1_U4 ( .A1(
        my_filter_delay_line_delay_chain_1_n51), .A2(
        my_filter_delay_line_delay_chain_1_n50), .ZN(
        my_filter_delay_line_delay_chain_1_n94) );
  BUF_X1 my_filter_delay_line_delay_chain_1_U3 ( .A(my_filter_delay_line_n11), 
        .Z(my_filter_delay_line_delay_chain_1_n51) );
  DFFR_X1 my_filter_delay_line_delay_chain_1_q_reg_0_ ( .D(
        my_filter_delay_line_delay_chain_1_n52), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_1_n51), .Q(
        my_filter_q_reg_chain_2__0_), .QN(
        my_filter_delay_line_delay_chain_1_n79) );
  DFFR_X1 my_filter_delay_line_delay_chain_1_q_reg_1_ ( .D(
        my_filter_delay_line_delay_chain_1_n53), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_1_n51), .Q(
        my_filter_q_reg_chain_2__1_), .QN(
        my_filter_delay_line_delay_chain_1_n78) );
  DFFR_X1 my_filter_delay_line_delay_chain_1_q_reg_2_ ( .D(
        my_filter_delay_line_delay_chain_1_n54), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_1_n51), .Q(
        my_filter_q_reg_chain_2__2_), .QN(
        my_filter_delay_line_delay_chain_1_n77) );
  DFFR_X1 my_filter_delay_line_delay_chain_1_q_reg_3_ ( .D(
        my_filter_delay_line_delay_chain_1_n55), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_1_n51), .Q(
        my_filter_q_reg_chain_2__3_), .QN(
        my_filter_delay_line_delay_chain_1_n76) );
  DFFR_X1 my_filter_delay_line_delay_chain_1_q_reg_4_ ( .D(
        my_filter_delay_line_delay_chain_1_n56), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_1_n51), .Q(
        my_filter_q_reg_chain_2__4_), .QN(
        my_filter_delay_line_delay_chain_1_n75) );
  DFFR_X1 my_filter_delay_line_delay_chain_1_q_reg_5_ ( .D(
        my_filter_delay_line_delay_chain_1_n57), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_1_n51), .Q(
        my_filter_q_reg_chain_2__5_), .QN(
        my_filter_delay_line_delay_chain_1_n74) );
  DFFR_X1 my_filter_delay_line_delay_chain_1_q_reg_6_ ( .D(
        my_filter_delay_line_delay_chain_1_n58), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_1_n51), .Q(
        my_filter_q_reg_chain_2__6_), .QN(
        my_filter_delay_line_delay_chain_1_n73) );
  DFFR_X1 my_filter_delay_line_delay_chain_1_q_reg_7_ ( .D(
        my_filter_delay_line_delay_chain_1_n59), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_1_n51), .Q(
        my_filter_q_reg_chain_2__7_), .QN(
        my_filter_delay_line_delay_chain_1_n72) );
  DFFR_X1 my_filter_delay_line_delay_chain_1_q_reg_8_ ( .D(
        my_filter_delay_line_delay_chain_1_n60), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_1_n51), .Q(
        my_filter_q_reg_chain_2__8_), .QN(
        my_filter_delay_line_delay_chain_1_n71) );
  DFFR_X1 my_filter_delay_line_delay_chain_1_q_reg_9_ ( .D(
        my_filter_delay_line_delay_chain_1_n61), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_1_n51), .Q(
        my_filter_q_reg_chain_2__9_), .QN(
        my_filter_delay_line_delay_chain_1_n70) );
  DFFR_X1 my_filter_delay_line_delay_chain_1_q_reg_10_ ( .D(
        my_filter_delay_line_delay_chain_1_n62), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_1_n51), .Q(
        my_filter_q_reg_chain_2__10_), .QN(
        my_filter_delay_line_delay_chain_1_n69) );
  DFFR_X1 my_filter_delay_line_delay_chain_1_q_reg_11_ ( .D(
        my_filter_delay_line_delay_chain_1_n63), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_1_n51), .Q(
        my_filter_q_reg_chain_2__11_), .QN(
        my_filter_delay_line_delay_chain_1_n68) );
  DFFR_X1 my_filter_delay_line_delay_chain_1_q_reg_12_ ( .D(
        my_filter_delay_line_delay_chain_1_n64), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_1_n51), .Q(
        my_filter_q_reg_chain_2__12_), .QN(
        my_filter_delay_line_delay_chain_1_n67) );
  DFFR_X1 my_filter_delay_line_delay_chain_1_q_reg_13_ ( .D(
        my_filter_delay_line_delay_chain_1_n65), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_1_n51), .Q(
        my_filter_q_reg_chain_2__13_), .QN(
        my_filter_delay_line_delay_chain_1_n66) );
  INV_X1 my_filter_delay_line_delay_chain_2_U35 ( .A(
        my_filter_delay_line_delay_chain_2_n50), .ZN(
        my_filter_delay_line_delay_chain_2_n49) );
  NAND2_X1 my_filter_delay_line_delay_chain_2_U34 ( .A1(
        my_filter_delay_line_delay_chain_2_n49), .A2(
        my_filter_q_reg_chain_2__13_), .ZN(
        my_filter_delay_line_delay_chain_2_n93) );
  OAI21_X1 my_filter_delay_line_delay_chain_2_U33 ( .B1(
        my_filter_delay_line_delay_chain_2_n94), .B2(
        my_filter_delay_line_delay_chain_2_n66), .A(
        my_filter_delay_line_delay_chain_2_n93), .ZN(
        my_filter_delay_line_delay_chain_2_n65) );
  NAND2_X1 my_filter_delay_line_delay_chain_2_U32 ( .A1(
        my_filter_q_reg_chain_2__12_), .A2(
        my_filter_delay_line_delay_chain_2_n49), .ZN(
        my_filter_delay_line_delay_chain_2_n92) );
  OAI21_X1 my_filter_delay_line_delay_chain_2_U31 ( .B1(
        my_filter_delay_line_delay_chain_2_n94), .B2(
        my_filter_delay_line_delay_chain_2_n67), .A(
        my_filter_delay_line_delay_chain_2_n92), .ZN(
        my_filter_delay_line_delay_chain_2_n64) );
  NAND2_X1 my_filter_delay_line_delay_chain_2_U30 ( .A1(
        my_filter_q_reg_chain_2__11_), .A2(
        my_filter_delay_line_delay_chain_2_n48), .ZN(
        my_filter_delay_line_delay_chain_2_n91) );
  OAI21_X1 my_filter_delay_line_delay_chain_2_U29 ( .B1(
        my_filter_delay_line_delay_chain_2_n94), .B2(
        my_filter_delay_line_delay_chain_2_n68), .A(
        my_filter_delay_line_delay_chain_2_n91), .ZN(
        my_filter_delay_line_delay_chain_2_n63) );
  NAND2_X1 my_filter_delay_line_delay_chain_2_U28 ( .A1(
        my_filter_q_reg_chain_2__10_), .A2(
        my_filter_delay_line_delay_chain_2_n48), .ZN(
        my_filter_delay_line_delay_chain_2_n90) );
  OAI21_X1 my_filter_delay_line_delay_chain_2_U27 ( .B1(
        my_filter_delay_line_delay_chain_2_n94), .B2(
        my_filter_delay_line_delay_chain_2_n69), .A(
        my_filter_delay_line_delay_chain_2_n90), .ZN(
        my_filter_delay_line_delay_chain_2_n62) );
  NAND2_X1 my_filter_delay_line_delay_chain_2_U26 ( .A1(
        my_filter_q_reg_chain_2__9_), .A2(
        my_filter_delay_line_delay_chain_2_n48), .ZN(
        my_filter_delay_line_delay_chain_2_n89) );
  OAI21_X1 my_filter_delay_line_delay_chain_2_U25 ( .B1(
        my_filter_delay_line_delay_chain_2_n94), .B2(
        my_filter_delay_line_delay_chain_2_n70), .A(
        my_filter_delay_line_delay_chain_2_n89), .ZN(
        my_filter_delay_line_delay_chain_2_n61) );
  NAND2_X1 my_filter_delay_line_delay_chain_2_U24 ( .A1(
        my_filter_q_reg_chain_2__8_), .A2(
        my_filter_delay_line_delay_chain_2_n48), .ZN(
        my_filter_delay_line_delay_chain_2_n88) );
  OAI21_X1 my_filter_delay_line_delay_chain_2_U23 ( .B1(
        my_filter_delay_line_delay_chain_2_n94), .B2(
        my_filter_delay_line_delay_chain_2_n71), .A(
        my_filter_delay_line_delay_chain_2_n88), .ZN(
        my_filter_delay_line_delay_chain_2_n60) );
  NAND2_X1 my_filter_delay_line_delay_chain_2_U22 ( .A1(
        my_filter_q_reg_chain_2__7_), .A2(
        my_filter_delay_line_delay_chain_2_n48), .ZN(
        my_filter_delay_line_delay_chain_2_n87) );
  OAI21_X1 my_filter_delay_line_delay_chain_2_U21 ( .B1(
        my_filter_delay_line_delay_chain_2_n94), .B2(
        my_filter_delay_line_delay_chain_2_n72), .A(
        my_filter_delay_line_delay_chain_2_n87), .ZN(
        my_filter_delay_line_delay_chain_2_n59) );
  NAND2_X1 my_filter_delay_line_delay_chain_2_U20 ( .A1(
        my_filter_q_reg_chain_2__6_), .A2(
        my_filter_delay_line_delay_chain_2_n48), .ZN(
        my_filter_delay_line_delay_chain_2_n86) );
  OAI21_X1 my_filter_delay_line_delay_chain_2_U19 ( .B1(
        my_filter_delay_line_delay_chain_2_n94), .B2(
        my_filter_delay_line_delay_chain_2_n73), .A(
        my_filter_delay_line_delay_chain_2_n86), .ZN(
        my_filter_delay_line_delay_chain_2_n58) );
  NAND2_X1 my_filter_delay_line_delay_chain_2_U18 ( .A1(
        my_filter_q_reg_chain_2__5_), .A2(
        my_filter_delay_line_delay_chain_2_n48), .ZN(
        my_filter_delay_line_delay_chain_2_n85) );
  OAI21_X1 my_filter_delay_line_delay_chain_2_U17 ( .B1(
        my_filter_delay_line_delay_chain_2_n94), .B2(
        my_filter_delay_line_delay_chain_2_n74), .A(
        my_filter_delay_line_delay_chain_2_n85), .ZN(
        my_filter_delay_line_delay_chain_2_n57) );
  NAND2_X1 my_filter_delay_line_delay_chain_2_U16 ( .A1(
        my_filter_q_reg_chain_2__4_), .A2(
        my_filter_delay_line_delay_chain_2_n48), .ZN(
        my_filter_delay_line_delay_chain_2_n84) );
  OAI21_X1 my_filter_delay_line_delay_chain_2_U15 ( .B1(
        my_filter_delay_line_delay_chain_2_n94), .B2(
        my_filter_delay_line_delay_chain_2_n75), .A(
        my_filter_delay_line_delay_chain_2_n84), .ZN(
        my_filter_delay_line_delay_chain_2_n56) );
  NAND2_X1 my_filter_delay_line_delay_chain_2_U14 ( .A1(
        my_filter_q_reg_chain_2__3_), .A2(
        my_filter_delay_line_delay_chain_2_n48), .ZN(
        my_filter_delay_line_delay_chain_2_n83) );
  OAI21_X1 my_filter_delay_line_delay_chain_2_U13 ( .B1(
        my_filter_delay_line_delay_chain_2_n94), .B2(
        my_filter_delay_line_delay_chain_2_n76), .A(
        my_filter_delay_line_delay_chain_2_n83), .ZN(
        my_filter_delay_line_delay_chain_2_n55) );
  NAND2_X1 my_filter_delay_line_delay_chain_2_U12 ( .A1(
        my_filter_q_reg_chain_2__2_), .A2(
        my_filter_delay_line_delay_chain_2_n48), .ZN(
        my_filter_delay_line_delay_chain_2_n82) );
  OAI21_X1 my_filter_delay_line_delay_chain_2_U11 ( .B1(
        my_filter_delay_line_delay_chain_2_n94), .B2(
        my_filter_delay_line_delay_chain_2_n77), .A(
        my_filter_delay_line_delay_chain_2_n82), .ZN(
        my_filter_delay_line_delay_chain_2_n54) );
  NAND2_X1 my_filter_delay_line_delay_chain_2_U10 ( .A1(
        my_filter_q_reg_chain_2__1_), .A2(
        my_filter_delay_line_delay_chain_2_n48), .ZN(
        my_filter_delay_line_delay_chain_2_n81) );
  OAI21_X1 my_filter_delay_line_delay_chain_2_U9 ( .B1(
        my_filter_delay_line_delay_chain_2_n94), .B2(
        my_filter_delay_line_delay_chain_2_n78), .A(
        my_filter_delay_line_delay_chain_2_n81), .ZN(
        my_filter_delay_line_delay_chain_2_n53) );
  NAND2_X1 my_filter_delay_line_delay_chain_2_U8 ( .A1(
        my_filter_q_reg_chain_2__0_), .A2(
        my_filter_delay_line_delay_chain_2_n48), .ZN(
        my_filter_delay_line_delay_chain_2_n80) );
  OAI21_X1 my_filter_delay_line_delay_chain_2_U7 ( .B1(
        my_filter_delay_line_delay_chain_2_n94), .B2(
        my_filter_delay_line_delay_chain_2_n79), .A(
        my_filter_delay_line_delay_chain_2_n80), .ZN(
        my_filter_delay_line_delay_chain_2_n52) );
  INV_X1 my_filter_delay_line_delay_chain_2_U6 ( .A(my_filter_delay_line_n8), 
        .ZN(my_filter_delay_line_delay_chain_2_n50) );
  INV_X1 my_filter_delay_line_delay_chain_2_U5 ( .A(
        my_filter_delay_line_delay_chain_2_n50), .ZN(
        my_filter_delay_line_delay_chain_2_n48) );
  NAND2_X1 my_filter_delay_line_delay_chain_2_U4 ( .A1(
        my_filter_delay_line_delay_chain_2_n51), .A2(
        my_filter_delay_line_delay_chain_2_n50), .ZN(
        my_filter_delay_line_delay_chain_2_n94) );
  BUF_X1 my_filter_delay_line_delay_chain_2_U3 ( .A(my_filter_delay_line_n11), 
        .Z(my_filter_delay_line_delay_chain_2_n51) );
  DFFR_X1 my_filter_delay_line_delay_chain_2_q_reg_0_ ( .D(
        my_filter_delay_line_delay_chain_2_n52), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_2_n51), .Q(
        my_filter_q_reg_chain_3__0_), .QN(
        my_filter_delay_line_delay_chain_2_n79) );
  DFFR_X1 my_filter_delay_line_delay_chain_2_q_reg_1_ ( .D(
        my_filter_delay_line_delay_chain_2_n53), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_2_n51), .Q(
        my_filter_q_reg_chain_3__1_), .QN(
        my_filter_delay_line_delay_chain_2_n78) );
  DFFR_X1 my_filter_delay_line_delay_chain_2_q_reg_2_ ( .D(
        my_filter_delay_line_delay_chain_2_n54), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_2_n51), .Q(
        my_filter_q_reg_chain_3__2_), .QN(
        my_filter_delay_line_delay_chain_2_n77) );
  DFFR_X1 my_filter_delay_line_delay_chain_2_q_reg_3_ ( .D(
        my_filter_delay_line_delay_chain_2_n55), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_2_n51), .Q(
        my_filter_q_reg_chain_3__3_), .QN(
        my_filter_delay_line_delay_chain_2_n76) );
  DFFR_X1 my_filter_delay_line_delay_chain_2_q_reg_4_ ( .D(
        my_filter_delay_line_delay_chain_2_n56), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_2_n51), .Q(
        my_filter_q_reg_chain_3__4_), .QN(
        my_filter_delay_line_delay_chain_2_n75) );
  DFFR_X1 my_filter_delay_line_delay_chain_2_q_reg_5_ ( .D(
        my_filter_delay_line_delay_chain_2_n57), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_2_n51), .Q(
        my_filter_q_reg_chain_3__5_), .QN(
        my_filter_delay_line_delay_chain_2_n74) );
  DFFR_X1 my_filter_delay_line_delay_chain_2_q_reg_6_ ( .D(
        my_filter_delay_line_delay_chain_2_n58), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_2_n51), .Q(
        my_filter_q_reg_chain_3__6_), .QN(
        my_filter_delay_line_delay_chain_2_n73) );
  DFFR_X1 my_filter_delay_line_delay_chain_2_q_reg_7_ ( .D(
        my_filter_delay_line_delay_chain_2_n59), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_2_n51), .Q(
        my_filter_q_reg_chain_3__7_), .QN(
        my_filter_delay_line_delay_chain_2_n72) );
  DFFR_X1 my_filter_delay_line_delay_chain_2_q_reg_8_ ( .D(
        my_filter_delay_line_delay_chain_2_n60), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_2_n51), .Q(
        my_filter_q_reg_chain_3__8_), .QN(
        my_filter_delay_line_delay_chain_2_n71) );
  DFFR_X1 my_filter_delay_line_delay_chain_2_q_reg_9_ ( .D(
        my_filter_delay_line_delay_chain_2_n61), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_2_n51), .Q(
        my_filter_q_reg_chain_3__9_), .QN(
        my_filter_delay_line_delay_chain_2_n70) );
  DFFR_X1 my_filter_delay_line_delay_chain_2_q_reg_10_ ( .D(
        my_filter_delay_line_delay_chain_2_n62), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_2_n51), .Q(
        my_filter_q_reg_chain_3__10_), .QN(
        my_filter_delay_line_delay_chain_2_n69) );
  DFFR_X1 my_filter_delay_line_delay_chain_2_q_reg_11_ ( .D(
        my_filter_delay_line_delay_chain_2_n63), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_2_n51), .Q(
        my_filter_q_reg_chain_3__11_), .QN(
        my_filter_delay_line_delay_chain_2_n68) );
  DFFR_X1 my_filter_delay_line_delay_chain_2_q_reg_12_ ( .D(
        my_filter_delay_line_delay_chain_2_n64), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_2_n51), .Q(
        my_filter_q_reg_chain_3__12_), .QN(
        my_filter_delay_line_delay_chain_2_n67) );
  DFFR_X1 my_filter_delay_line_delay_chain_2_q_reg_13_ ( .D(
        my_filter_delay_line_delay_chain_2_n65), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_2_n51), .Q(
        my_filter_q_reg_chain_3__13_), .QN(
        my_filter_delay_line_delay_chain_2_n66) );
  INV_X1 my_filter_delay_line_delay_chain_3_U35 ( .A(
        my_filter_delay_line_delay_chain_3_n50), .ZN(
        my_filter_delay_line_delay_chain_3_n49) );
  NAND2_X1 my_filter_delay_line_delay_chain_3_U34 ( .A1(
        my_filter_delay_line_delay_chain_3_n49), .A2(
        my_filter_q_reg_chain_3__13_), .ZN(
        my_filter_delay_line_delay_chain_3_n93) );
  OAI21_X1 my_filter_delay_line_delay_chain_3_U33 ( .B1(
        my_filter_delay_line_delay_chain_3_n94), .B2(
        my_filter_delay_line_delay_chain_3_n66), .A(
        my_filter_delay_line_delay_chain_3_n93), .ZN(
        my_filter_delay_line_delay_chain_3_n65) );
  NAND2_X1 my_filter_delay_line_delay_chain_3_U32 ( .A1(
        my_filter_q_reg_chain_3__12_), .A2(
        my_filter_delay_line_delay_chain_3_n49), .ZN(
        my_filter_delay_line_delay_chain_3_n92) );
  OAI21_X1 my_filter_delay_line_delay_chain_3_U31 ( .B1(
        my_filter_delay_line_delay_chain_3_n94), .B2(
        my_filter_delay_line_delay_chain_3_n67), .A(
        my_filter_delay_line_delay_chain_3_n92), .ZN(
        my_filter_delay_line_delay_chain_3_n64) );
  NAND2_X1 my_filter_delay_line_delay_chain_3_U30 ( .A1(
        my_filter_q_reg_chain_3__11_), .A2(
        my_filter_delay_line_delay_chain_3_n48), .ZN(
        my_filter_delay_line_delay_chain_3_n91) );
  OAI21_X1 my_filter_delay_line_delay_chain_3_U29 ( .B1(
        my_filter_delay_line_delay_chain_3_n94), .B2(
        my_filter_delay_line_delay_chain_3_n68), .A(
        my_filter_delay_line_delay_chain_3_n91), .ZN(
        my_filter_delay_line_delay_chain_3_n63) );
  NAND2_X1 my_filter_delay_line_delay_chain_3_U28 ( .A1(
        my_filter_q_reg_chain_3__10_), .A2(
        my_filter_delay_line_delay_chain_3_n48), .ZN(
        my_filter_delay_line_delay_chain_3_n90) );
  OAI21_X1 my_filter_delay_line_delay_chain_3_U27 ( .B1(
        my_filter_delay_line_delay_chain_3_n94), .B2(
        my_filter_delay_line_delay_chain_3_n69), .A(
        my_filter_delay_line_delay_chain_3_n90), .ZN(
        my_filter_delay_line_delay_chain_3_n62) );
  NAND2_X1 my_filter_delay_line_delay_chain_3_U26 ( .A1(
        my_filter_q_reg_chain_3__9_), .A2(
        my_filter_delay_line_delay_chain_3_n48), .ZN(
        my_filter_delay_line_delay_chain_3_n89) );
  OAI21_X1 my_filter_delay_line_delay_chain_3_U25 ( .B1(
        my_filter_delay_line_delay_chain_3_n94), .B2(
        my_filter_delay_line_delay_chain_3_n70), .A(
        my_filter_delay_line_delay_chain_3_n89), .ZN(
        my_filter_delay_line_delay_chain_3_n61) );
  NAND2_X1 my_filter_delay_line_delay_chain_3_U24 ( .A1(
        my_filter_q_reg_chain_3__8_), .A2(
        my_filter_delay_line_delay_chain_3_n48), .ZN(
        my_filter_delay_line_delay_chain_3_n88) );
  OAI21_X1 my_filter_delay_line_delay_chain_3_U23 ( .B1(
        my_filter_delay_line_delay_chain_3_n94), .B2(
        my_filter_delay_line_delay_chain_3_n71), .A(
        my_filter_delay_line_delay_chain_3_n88), .ZN(
        my_filter_delay_line_delay_chain_3_n60) );
  NAND2_X1 my_filter_delay_line_delay_chain_3_U22 ( .A1(
        my_filter_q_reg_chain_3__7_), .A2(
        my_filter_delay_line_delay_chain_3_n48), .ZN(
        my_filter_delay_line_delay_chain_3_n87) );
  OAI21_X1 my_filter_delay_line_delay_chain_3_U21 ( .B1(
        my_filter_delay_line_delay_chain_3_n94), .B2(
        my_filter_delay_line_delay_chain_3_n72), .A(
        my_filter_delay_line_delay_chain_3_n87), .ZN(
        my_filter_delay_line_delay_chain_3_n59) );
  NAND2_X1 my_filter_delay_line_delay_chain_3_U20 ( .A1(
        my_filter_q_reg_chain_3__6_), .A2(
        my_filter_delay_line_delay_chain_3_n48), .ZN(
        my_filter_delay_line_delay_chain_3_n86) );
  OAI21_X1 my_filter_delay_line_delay_chain_3_U19 ( .B1(
        my_filter_delay_line_delay_chain_3_n94), .B2(
        my_filter_delay_line_delay_chain_3_n73), .A(
        my_filter_delay_line_delay_chain_3_n86), .ZN(
        my_filter_delay_line_delay_chain_3_n58) );
  NAND2_X1 my_filter_delay_line_delay_chain_3_U18 ( .A1(
        my_filter_q_reg_chain_3__5_), .A2(
        my_filter_delay_line_delay_chain_3_n48), .ZN(
        my_filter_delay_line_delay_chain_3_n85) );
  OAI21_X1 my_filter_delay_line_delay_chain_3_U17 ( .B1(
        my_filter_delay_line_delay_chain_3_n94), .B2(
        my_filter_delay_line_delay_chain_3_n74), .A(
        my_filter_delay_line_delay_chain_3_n85), .ZN(
        my_filter_delay_line_delay_chain_3_n57) );
  NAND2_X1 my_filter_delay_line_delay_chain_3_U16 ( .A1(
        my_filter_q_reg_chain_3__4_), .A2(
        my_filter_delay_line_delay_chain_3_n48), .ZN(
        my_filter_delay_line_delay_chain_3_n84) );
  OAI21_X1 my_filter_delay_line_delay_chain_3_U15 ( .B1(
        my_filter_delay_line_delay_chain_3_n94), .B2(
        my_filter_delay_line_delay_chain_3_n75), .A(
        my_filter_delay_line_delay_chain_3_n84), .ZN(
        my_filter_delay_line_delay_chain_3_n56) );
  NAND2_X1 my_filter_delay_line_delay_chain_3_U14 ( .A1(
        my_filter_q_reg_chain_3__3_), .A2(
        my_filter_delay_line_delay_chain_3_n48), .ZN(
        my_filter_delay_line_delay_chain_3_n83) );
  OAI21_X1 my_filter_delay_line_delay_chain_3_U13 ( .B1(
        my_filter_delay_line_delay_chain_3_n94), .B2(
        my_filter_delay_line_delay_chain_3_n76), .A(
        my_filter_delay_line_delay_chain_3_n83), .ZN(
        my_filter_delay_line_delay_chain_3_n55) );
  NAND2_X1 my_filter_delay_line_delay_chain_3_U12 ( .A1(
        my_filter_q_reg_chain_3__2_), .A2(
        my_filter_delay_line_delay_chain_3_n48), .ZN(
        my_filter_delay_line_delay_chain_3_n82) );
  OAI21_X1 my_filter_delay_line_delay_chain_3_U11 ( .B1(
        my_filter_delay_line_delay_chain_3_n94), .B2(
        my_filter_delay_line_delay_chain_3_n77), .A(
        my_filter_delay_line_delay_chain_3_n82), .ZN(
        my_filter_delay_line_delay_chain_3_n54) );
  NAND2_X1 my_filter_delay_line_delay_chain_3_U10 ( .A1(
        my_filter_q_reg_chain_3__1_), .A2(
        my_filter_delay_line_delay_chain_3_n48), .ZN(
        my_filter_delay_line_delay_chain_3_n81) );
  OAI21_X1 my_filter_delay_line_delay_chain_3_U9 ( .B1(
        my_filter_delay_line_delay_chain_3_n94), .B2(
        my_filter_delay_line_delay_chain_3_n78), .A(
        my_filter_delay_line_delay_chain_3_n81), .ZN(
        my_filter_delay_line_delay_chain_3_n53) );
  NAND2_X1 my_filter_delay_line_delay_chain_3_U8 ( .A1(
        my_filter_q_reg_chain_3__0_), .A2(
        my_filter_delay_line_delay_chain_3_n48), .ZN(
        my_filter_delay_line_delay_chain_3_n80) );
  OAI21_X1 my_filter_delay_line_delay_chain_3_U7 ( .B1(
        my_filter_delay_line_delay_chain_3_n94), .B2(
        my_filter_delay_line_delay_chain_3_n79), .A(
        my_filter_delay_line_delay_chain_3_n80), .ZN(
        my_filter_delay_line_delay_chain_3_n52) );
  INV_X1 my_filter_delay_line_delay_chain_3_U6 ( .A(my_filter_delay_line_n8), 
        .ZN(my_filter_delay_line_delay_chain_3_n50) );
  INV_X1 my_filter_delay_line_delay_chain_3_U5 ( .A(
        my_filter_delay_line_delay_chain_3_n50), .ZN(
        my_filter_delay_line_delay_chain_3_n48) );
  NAND2_X1 my_filter_delay_line_delay_chain_3_U4 ( .A1(
        my_filter_delay_line_delay_chain_3_n51), .A2(
        my_filter_delay_line_delay_chain_3_n50), .ZN(
        my_filter_delay_line_delay_chain_3_n94) );
  BUF_X1 my_filter_delay_line_delay_chain_3_U3 ( .A(my_filter_delay_line_n12), 
        .Z(my_filter_delay_line_delay_chain_3_n51) );
  DFFR_X1 my_filter_delay_line_delay_chain_3_q_reg_0_ ( .D(
        my_filter_delay_line_delay_chain_3_n52), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_3_n51), .Q(
        my_filter_q_reg_chain_4__0_), .QN(
        my_filter_delay_line_delay_chain_3_n79) );
  DFFR_X1 my_filter_delay_line_delay_chain_3_q_reg_1_ ( .D(
        my_filter_delay_line_delay_chain_3_n53), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_3_n51), .Q(
        my_filter_q_reg_chain_4__1_), .QN(
        my_filter_delay_line_delay_chain_3_n78) );
  DFFR_X1 my_filter_delay_line_delay_chain_3_q_reg_2_ ( .D(
        my_filter_delay_line_delay_chain_3_n54), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_3_n51), .Q(
        my_filter_q_reg_chain_4__2_), .QN(
        my_filter_delay_line_delay_chain_3_n77) );
  DFFR_X1 my_filter_delay_line_delay_chain_3_q_reg_3_ ( .D(
        my_filter_delay_line_delay_chain_3_n55), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_3_n51), .Q(
        my_filter_q_reg_chain_4__3_), .QN(
        my_filter_delay_line_delay_chain_3_n76) );
  DFFR_X1 my_filter_delay_line_delay_chain_3_q_reg_4_ ( .D(
        my_filter_delay_line_delay_chain_3_n56), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_3_n51), .Q(
        my_filter_q_reg_chain_4__4_), .QN(
        my_filter_delay_line_delay_chain_3_n75) );
  DFFR_X1 my_filter_delay_line_delay_chain_3_q_reg_5_ ( .D(
        my_filter_delay_line_delay_chain_3_n57), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_3_n51), .Q(
        my_filter_q_reg_chain_4__5_), .QN(
        my_filter_delay_line_delay_chain_3_n74) );
  DFFR_X1 my_filter_delay_line_delay_chain_3_q_reg_6_ ( .D(
        my_filter_delay_line_delay_chain_3_n58), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_3_n51), .Q(
        my_filter_q_reg_chain_4__6_), .QN(
        my_filter_delay_line_delay_chain_3_n73) );
  DFFR_X1 my_filter_delay_line_delay_chain_3_q_reg_7_ ( .D(
        my_filter_delay_line_delay_chain_3_n59), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_3_n51), .Q(
        my_filter_q_reg_chain_4__7_), .QN(
        my_filter_delay_line_delay_chain_3_n72) );
  DFFR_X1 my_filter_delay_line_delay_chain_3_q_reg_8_ ( .D(
        my_filter_delay_line_delay_chain_3_n60), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_3_n51), .Q(
        my_filter_q_reg_chain_4__8_), .QN(
        my_filter_delay_line_delay_chain_3_n71) );
  DFFR_X1 my_filter_delay_line_delay_chain_3_q_reg_9_ ( .D(
        my_filter_delay_line_delay_chain_3_n61), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_3_n51), .Q(
        my_filter_q_reg_chain_4__9_), .QN(
        my_filter_delay_line_delay_chain_3_n70) );
  DFFR_X1 my_filter_delay_line_delay_chain_3_q_reg_10_ ( .D(
        my_filter_delay_line_delay_chain_3_n62), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_3_n51), .Q(
        my_filter_q_reg_chain_4__10_), .QN(
        my_filter_delay_line_delay_chain_3_n69) );
  DFFR_X1 my_filter_delay_line_delay_chain_3_q_reg_11_ ( .D(
        my_filter_delay_line_delay_chain_3_n63), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_3_n51), .Q(
        my_filter_q_reg_chain_4__11_), .QN(
        my_filter_delay_line_delay_chain_3_n68) );
  DFFR_X1 my_filter_delay_line_delay_chain_3_q_reg_12_ ( .D(
        my_filter_delay_line_delay_chain_3_n64), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_3_n51), .Q(
        my_filter_q_reg_chain_4__12_), .QN(
        my_filter_delay_line_delay_chain_3_n67) );
  DFFR_X1 my_filter_delay_line_delay_chain_3_q_reg_13_ ( .D(
        my_filter_delay_line_delay_chain_3_n65), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_3_n51), .Q(
        my_filter_q_reg_chain_4__13_), .QN(
        my_filter_delay_line_delay_chain_3_n66) );
  INV_X1 my_filter_delay_line_delay_chain_4_U35 ( .A(
        my_filter_delay_line_delay_chain_4_n50), .ZN(
        my_filter_delay_line_delay_chain_4_n49) );
  NAND2_X1 my_filter_delay_line_delay_chain_4_U34 ( .A1(
        my_filter_delay_line_delay_chain_4_n49), .A2(
        my_filter_q_reg_chain_4__13_), .ZN(
        my_filter_delay_line_delay_chain_4_n93) );
  OAI21_X1 my_filter_delay_line_delay_chain_4_U33 ( .B1(
        my_filter_delay_line_delay_chain_4_n94), .B2(
        my_filter_delay_line_delay_chain_4_n66), .A(
        my_filter_delay_line_delay_chain_4_n93), .ZN(
        my_filter_delay_line_delay_chain_4_n65) );
  NAND2_X1 my_filter_delay_line_delay_chain_4_U32 ( .A1(
        my_filter_q_reg_chain_4__12_), .A2(
        my_filter_delay_line_delay_chain_4_n49), .ZN(
        my_filter_delay_line_delay_chain_4_n92) );
  OAI21_X1 my_filter_delay_line_delay_chain_4_U31 ( .B1(
        my_filter_delay_line_delay_chain_4_n94), .B2(
        my_filter_delay_line_delay_chain_4_n67), .A(
        my_filter_delay_line_delay_chain_4_n92), .ZN(
        my_filter_delay_line_delay_chain_4_n64) );
  NAND2_X1 my_filter_delay_line_delay_chain_4_U30 ( .A1(
        my_filter_q_reg_chain_4__11_), .A2(
        my_filter_delay_line_delay_chain_4_n48), .ZN(
        my_filter_delay_line_delay_chain_4_n91) );
  OAI21_X1 my_filter_delay_line_delay_chain_4_U29 ( .B1(
        my_filter_delay_line_delay_chain_4_n94), .B2(
        my_filter_delay_line_delay_chain_4_n68), .A(
        my_filter_delay_line_delay_chain_4_n91), .ZN(
        my_filter_delay_line_delay_chain_4_n63) );
  NAND2_X1 my_filter_delay_line_delay_chain_4_U28 ( .A1(
        my_filter_q_reg_chain_4__10_), .A2(
        my_filter_delay_line_delay_chain_4_n48), .ZN(
        my_filter_delay_line_delay_chain_4_n90) );
  OAI21_X1 my_filter_delay_line_delay_chain_4_U27 ( .B1(
        my_filter_delay_line_delay_chain_4_n94), .B2(
        my_filter_delay_line_delay_chain_4_n69), .A(
        my_filter_delay_line_delay_chain_4_n90), .ZN(
        my_filter_delay_line_delay_chain_4_n62) );
  NAND2_X1 my_filter_delay_line_delay_chain_4_U26 ( .A1(
        my_filter_q_reg_chain_4__9_), .A2(
        my_filter_delay_line_delay_chain_4_n48), .ZN(
        my_filter_delay_line_delay_chain_4_n89) );
  OAI21_X1 my_filter_delay_line_delay_chain_4_U25 ( .B1(
        my_filter_delay_line_delay_chain_4_n94), .B2(
        my_filter_delay_line_delay_chain_4_n70), .A(
        my_filter_delay_line_delay_chain_4_n89), .ZN(
        my_filter_delay_line_delay_chain_4_n61) );
  NAND2_X1 my_filter_delay_line_delay_chain_4_U24 ( .A1(
        my_filter_q_reg_chain_4__8_), .A2(
        my_filter_delay_line_delay_chain_4_n48), .ZN(
        my_filter_delay_line_delay_chain_4_n88) );
  OAI21_X1 my_filter_delay_line_delay_chain_4_U23 ( .B1(
        my_filter_delay_line_delay_chain_4_n94), .B2(
        my_filter_delay_line_delay_chain_4_n71), .A(
        my_filter_delay_line_delay_chain_4_n88), .ZN(
        my_filter_delay_line_delay_chain_4_n60) );
  NAND2_X1 my_filter_delay_line_delay_chain_4_U22 ( .A1(
        my_filter_q_reg_chain_4__7_), .A2(
        my_filter_delay_line_delay_chain_4_n48), .ZN(
        my_filter_delay_line_delay_chain_4_n87) );
  OAI21_X1 my_filter_delay_line_delay_chain_4_U21 ( .B1(
        my_filter_delay_line_delay_chain_4_n94), .B2(
        my_filter_delay_line_delay_chain_4_n72), .A(
        my_filter_delay_line_delay_chain_4_n87), .ZN(
        my_filter_delay_line_delay_chain_4_n59) );
  NAND2_X1 my_filter_delay_line_delay_chain_4_U20 ( .A1(
        my_filter_q_reg_chain_4__6_), .A2(
        my_filter_delay_line_delay_chain_4_n48), .ZN(
        my_filter_delay_line_delay_chain_4_n86) );
  OAI21_X1 my_filter_delay_line_delay_chain_4_U19 ( .B1(
        my_filter_delay_line_delay_chain_4_n94), .B2(
        my_filter_delay_line_delay_chain_4_n73), .A(
        my_filter_delay_line_delay_chain_4_n86), .ZN(
        my_filter_delay_line_delay_chain_4_n58) );
  NAND2_X1 my_filter_delay_line_delay_chain_4_U18 ( .A1(
        my_filter_q_reg_chain_4__5_), .A2(
        my_filter_delay_line_delay_chain_4_n48), .ZN(
        my_filter_delay_line_delay_chain_4_n85) );
  OAI21_X1 my_filter_delay_line_delay_chain_4_U17 ( .B1(
        my_filter_delay_line_delay_chain_4_n94), .B2(
        my_filter_delay_line_delay_chain_4_n74), .A(
        my_filter_delay_line_delay_chain_4_n85), .ZN(
        my_filter_delay_line_delay_chain_4_n57) );
  NAND2_X1 my_filter_delay_line_delay_chain_4_U16 ( .A1(
        my_filter_q_reg_chain_4__4_), .A2(
        my_filter_delay_line_delay_chain_4_n48), .ZN(
        my_filter_delay_line_delay_chain_4_n84) );
  OAI21_X1 my_filter_delay_line_delay_chain_4_U15 ( .B1(
        my_filter_delay_line_delay_chain_4_n94), .B2(
        my_filter_delay_line_delay_chain_4_n75), .A(
        my_filter_delay_line_delay_chain_4_n84), .ZN(
        my_filter_delay_line_delay_chain_4_n56) );
  NAND2_X1 my_filter_delay_line_delay_chain_4_U14 ( .A1(
        my_filter_q_reg_chain_4__3_), .A2(
        my_filter_delay_line_delay_chain_4_n48), .ZN(
        my_filter_delay_line_delay_chain_4_n83) );
  OAI21_X1 my_filter_delay_line_delay_chain_4_U13 ( .B1(
        my_filter_delay_line_delay_chain_4_n94), .B2(
        my_filter_delay_line_delay_chain_4_n76), .A(
        my_filter_delay_line_delay_chain_4_n83), .ZN(
        my_filter_delay_line_delay_chain_4_n55) );
  NAND2_X1 my_filter_delay_line_delay_chain_4_U12 ( .A1(
        my_filter_q_reg_chain_4__2_), .A2(
        my_filter_delay_line_delay_chain_4_n48), .ZN(
        my_filter_delay_line_delay_chain_4_n82) );
  OAI21_X1 my_filter_delay_line_delay_chain_4_U11 ( .B1(
        my_filter_delay_line_delay_chain_4_n94), .B2(
        my_filter_delay_line_delay_chain_4_n77), .A(
        my_filter_delay_line_delay_chain_4_n82), .ZN(
        my_filter_delay_line_delay_chain_4_n54) );
  NAND2_X1 my_filter_delay_line_delay_chain_4_U10 ( .A1(
        my_filter_q_reg_chain_4__1_), .A2(
        my_filter_delay_line_delay_chain_4_n48), .ZN(
        my_filter_delay_line_delay_chain_4_n81) );
  OAI21_X1 my_filter_delay_line_delay_chain_4_U9 ( .B1(
        my_filter_delay_line_delay_chain_4_n94), .B2(
        my_filter_delay_line_delay_chain_4_n78), .A(
        my_filter_delay_line_delay_chain_4_n81), .ZN(
        my_filter_delay_line_delay_chain_4_n53) );
  NAND2_X1 my_filter_delay_line_delay_chain_4_U8 ( .A1(
        my_filter_q_reg_chain_4__0_), .A2(
        my_filter_delay_line_delay_chain_4_n48), .ZN(
        my_filter_delay_line_delay_chain_4_n80) );
  OAI21_X1 my_filter_delay_line_delay_chain_4_U7 ( .B1(
        my_filter_delay_line_delay_chain_4_n94), .B2(
        my_filter_delay_line_delay_chain_4_n79), .A(
        my_filter_delay_line_delay_chain_4_n80), .ZN(
        my_filter_delay_line_delay_chain_4_n52) );
  INV_X1 my_filter_delay_line_delay_chain_4_U6 ( .A(my_filter_delay_line_n8), 
        .ZN(my_filter_delay_line_delay_chain_4_n50) );
  INV_X1 my_filter_delay_line_delay_chain_4_U5 ( .A(
        my_filter_delay_line_delay_chain_4_n50), .ZN(
        my_filter_delay_line_delay_chain_4_n48) );
  NAND2_X1 my_filter_delay_line_delay_chain_4_U4 ( .A1(
        my_filter_delay_line_delay_chain_4_n51), .A2(
        my_filter_delay_line_delay_chain_4_n50), .ZN(
        my_filter_delay_line_delay_chain_4_n94) );
  BUF_X1 my_filter_delay_line_delay_chain_4_U3 ( .A(my_filter_delay_line_n12), 
        .Z(my_filter_delay_line_delay_chain_4_n51) );
  DFFR_X1 my_filter_delay_line_delay_chain_4_q_reg_0_ ( .D(
        my_filter_delay_line_delay_chain_4_n52), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_4_n51), .Q(
        my_filter_q_reg_chain_5__0_), .QN(
        my_filter_delay_line_delay_chain_4_n79) );
  DFFR_X1 my_filter_delay_line_delay_chain_4_q_reg_1_ ( .D(
        my_filter_delay_line_delay_chain_4_n53), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_4_n51), .Q(
        my_filter_q_reg_chain_5__1_), .QN(
        my_filter_delay_line_delay_chain_4_n78) );
  DFFR_X1 my_filter_delay_line_delay_chain_4_q_reg_2_ ( .D(
        my_filter_delay_line_delay_chain_4_n54), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_4_n51), .Q(
        my_filter_q_reg_chain_5__2_), .QN(
        my_filter_delay_line_delay_chain_4_n77) );
  DFFR_X1 my_filter_delay_line_delay_chain_4_q_reg_3_ ( .D(
        my_filter_delay_line_delay_chain_4_n55), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_4_n51), .Q(
        my_filter_q_reg_chain_5__3_), .QN(
        my_filter_delay_line_delay_chain_4_n76) );
  DFFR_X1 my_filter_delay_line_delay_chain_4_q_reg_4_ ( .D(
        my_filter_delay_line_delay_chain_4_n56), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_4_n51), .Q(
        my_filter_q_reg_chain_5__4_), .QN(
        my_filter_delay_line_delay_chain_4_n75) );
  DFFR_X1 my_filter_delay_line_delay_chain_4_q_reg_5_ ( .D(
        my_filter_delay_line_delay_chain_4_n57), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_4_n51), .Q(
        my_filter_q_reg_chain_5__5_), .QN(
        my_filter_delay_line_delay_chain_4_n74) );
  DFFR_X1 my_filter_delay_line_delay_chain_4_q_reg_6_ ( .D(
        my_filter_delay_line_delay_chain_4_n58), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_4_n51), .Q(
        my_filter_q_reg_chain_5__6_), .QN(
        my_filter_delay_line_delay_chain_4_n73) );
  DFFR_X1 my_filter_delay_line_delay_chain_4_q_reg_7_ ( .D(
        my_filter_delay_line_delay_chain_4_n59), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_4_n51), .Q(
        my_filter_q_reg_chain_5__7_), .QN(
        my_filter_delay_line_delay_chain_4_n72) );
  DFFR_X1 my_filter_delay_line_delay_chain_4_q_reg_8_ ( .D(
        my_filter_delay_line_delay_chain_4_n60), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_4_n51), .Q(
        my_filter_q_reg_chain_5__8_), .QN(
        my_filter_delay_line_delay_chain_4_n71) );
  DFFR_X1 my_filter_delay_line_delay_chain_4_q_reg_9_ ( .D(
        my_filter_delay_line_delay_chain_4_n61), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_4_n51), .Q(
        my_filter_q_reg_chain_5__9_), .QN(
        my_filter_delay_line_delay_chain_4_n70) );
  DFFR_X1 my_filter_delay_line_delay_chain_4_q_reg_10_ ( .D(
        my_filter_delay_line_delay_chain_4_n62), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_4_n51), .Q(
        my_filter_q_reg_chain_5__10_), .QN(
        my_filter_delay_line_delay_chain_4_n69) );
  DFFR_X1 my_filter_delay_line_delay_chain_4_q_reg_11_ ( .D(
        my_filter_delay_line_delay_chain_4_n63), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_4_n51), .Q(
        my_filter_q_reg_chain_5__11_), .QN(
        my_filter_delay_line_delay_chain_4_n68) );
  DFFR_X1 my_filter_delay_line_delay_chain_4_q_reg_12_ ( .D(
        my_filter_delay_line_delay_chain_4_n64), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_4_n51), .Q(
        my_filter_q_reg_chain_5__12_), .QN(
        my_filter_delay_line_delay_chain_4_n67) );
  DFFR_X1 my_filter_delay_line_delay_chain_4_q_reg_13_ ( .D(
        my_filter_delay_line_delay_chain_4_n65), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_4_n51), .Q(
        my_filter_q_reg_chain_5__13_), .QN(
        my_filter_delay_line_delay_chain_4_n66) );
  INV_X1 my_filter_delay_line_delay_chain_5_U35 ( .A(
        my_filter_delay_line_delay_chain_5_n50), .ZN(
        my_filter_delay_line_delay_chain_5_n49) );
  NAND2_X1 my_filter_delay_line_delay_chain_5_U34 ( .A1(
        my_filter_delay_line_delay_chain_5_n49), .A2(
        my_filter_q_reg_chain_5__13_), .ZN(
        my_filter_delay_line_delay_chain_5_n93) );
  OAI21_X1 my_filter_delay_line_delay_chain_5_U33 ( .B1(
        my_filter_delay_line_delay_chain_5_n94), .B2(
        my_filter_delay_line_delay_chain_5_n66), .A(
        my_filter_delay_line_delay_chain_5_n93), .ZN(
        my_filter_delay_line_delay_chain_5_n65) );
  NAND2_X1 my_filter_delay_line_delay_chain_5_U32 ( .A1(
        my_filter_q_reg_chain_5__12_), .A2(
        my_filter_delay_line_delay_chain_5_n49), .ZN(
        my_filter_delay_line_delay_chain_5_n92) );
  OAI21_X1 my_filter_delay_line_delay_chain_5_U31 ( .B1(
        my_filter_delay_line_delay_chain_5_n94), .B2(
        my_filter_delay_line_delay_chain_5_n67), .A(
        my_filter_delay_line_delay_chain_5_n92), .ZN(
        my_filter_delay_line_delay_chain_5_n64) );
  NAND2_X1 my_filter_delay_line_delay_chain_5_U30 ( .A1(
        my_filter_q_reg_chain_5__11_), .A2(
        my_filter_delay_line_delay_chain_5_n48), .ZN(
        my_filter_delay_line_delay_chain_5_n91) );
  OAI21_X1 my_filter_delay_line_delay_chain_5_U29 ( .B1(
        my_filter_delay_line_delay_chain_5_n94), .B2(
        my_filter_delay_line_delay_chain_5_n68), .A(
        my_filter_delay_line_delay_chain_5_n91), .ZN(
        my_filter_delay_line_delay_chain_5_n63) );
  NAND2_X1 my_filter_delay_line_delay_chain_5_U28 ( .A1(
        my_filter_q_reg_chain_5__10_), .A2(
        my_filter_delay_line_delay_chain_5_n48), .ZN(
        my_filter_delay_line_delay_chain_5_n90) );
  OAI21_X1 my_filter_delay_line_delay_chain_5_U27 ( .B1(
        my_filter_delay_line_delay_chain_5_n94), .B2(
        my_filter_delay_line_delay_chain_5_n69), .A(
        my_filter_delay_line_delay_chain_5_n90), .ZN(
        my_filter_delay_line_delay_chain_5_n62) );
  NAND2_X1 my_filter_delay_line_delay_chain_5_U26 ( .A1(
        my_filter_q_reg_chain_5__9_), .A2(
        my_filter_delay_line_delay_chain_5_n48), .ZN(
        my_filter_delay_line_delay_chain_5_n89) );
  OAI21_X1 my_filter_delay_line_delay_chain_5_U25 ( .B1(
        my_filter_delay_line_delay_chain_5_n94), .B2(
        my_filter_delay_line_delay_chain_5_n70), .A(
        my_filter_delay_line_delay_chain_5_n89), .ZN(
        my_filter_delay_line_delay_chain_5_n61) );
  NAND2_X1 my_filter_delay_line_delay_chain_5_U24 ( .A1(
        my_filter_q_reg_chain_5__8_), .A2(
        my_filter_delay_line_delay_chain_5_n48), .ZN(
        my_filter_delay_line_delay_chain_5_n88) );
  OAI21_X1 my_filter_delay_line_delay_chain_5_U23 ( .B1(
        my_filter_delay_line_delay_chain_5_n94), .B2(
        my_filter_delay_line_delay_chain_5_n71), .A(
        my_filter_delay_line_delay_chain_5_n88), .ZN(
        my_filter_delay_line_delay_chain_5_n60) );
  NAND2_X1 my_filter_delay_line_delay_chain_5_U22 ( .A1(
        my_filter_q_reg_chain_5__7_), .A2(
        my_filter_delay_line_delay_chain_5_n48), .ZN(
        my_filter_delay_line_delay_chain_5_n87) );
  OAI21_X1 my_filter_delay_line_delay_chain_5_U21 ( .B1(
        my_filter_delay_line_delay_chain_5_n94), .B2(
        my_filter_delay_line_delay_chain_5_n72), .A(
        my_filter_delay_line_delay_chain_5_n87), .ZN(
        my_filter_delay_line_delay_chain_5_n59) );
  NAND2_X1 my_filter_delay_line_delay_chain_5_U20 ( .A1(
        my_filter_q_reg_chain_5__6_), .A2(
        my_filter_delay_line_delay_chain_5_n48), .ZN(
        my_filter_delay_line_delay_chain_5_n86) );
  OAI21_X1 my_filter_delay_line_delay_chain_5_U19 ( .B1(
        my_filter_delay_line_delay_chain_5_n94), .B2(
        my_filter_delay_line_delay_chain_5_n73), .A(
        my_filter_delay_line_delay_chain_5_n86), .ZN(
        my_filter_delay_line_delay_chain_5_n58) );
  NAND2_X1 my_filter_delay_line_delay_chain_5_U18 ( .A1(
        my_filter_q_reg_chain_5__5_), .A2(
        my_filter_delay_line_delay_chain_5_n48), .ZN(
        my_filter_delay_line_delay_chain_5_n85) );
  OAI21_X1 my_filter_delay_line_delay_chain_5_U17 ( .B1(
        my_filter_delay_line_delay_chain_5_n94), .B2(
        my_filter_delay_line_delay_chain_5_n74), .A(
        my_filter_delay_line_delay_chain_5_n85), .ZN(
        my_filter_delay_line_delay_chain_5_n57) );
  NAND2_X1 my_filter_delay_line_delay_chain_5_U16 ( .A1(
        my_filter_q_reg_chain_5__4_), .A2(
        my_filter_delay_line_delay_chain_5_n48), .ZN(
        my_filter_delay_line_delay_chain_5_n84) );
  OAI21_X1 my_filter_delay_line_delay_chain_5_U15 ( .B1(
        my_filter_delay_line_delay_chain_5_n94), .B2(
        my_filter_delay_line_delay_chain_5_n75), .A(
        my_filter_delay_line_delay_chain_5_n84), .ZN(
        my_filter_delay_line_delay_chain_5_n56) );
  NAND2_X1 my_filter_delay_line_delay_chain_5_U14 ( .A1(
        my_filter_q_reg_chain_5__3_), .A2(
        my_filter_delay_line_delay_chain_5_n48), .ZN(
        my_filter_delay_line_delay_chain_5_n83) );
  OAI21_X1 my_filter_delay_line_delay_chain_5_U13 ( .B1(
        my_filter_delay_line_delay_chain_5_n94), .B2(
        my_filter_delay_line_delay_chain_5_n76), .A(
        my_filter_delay_line_delay_chain_5_n83), .ZN(
        my_filter_delay_line_delay_chain_5_n55) );
  NAND2_X1 my_filter_delay_line_delay_chain_5_U12 ( .A1(
        my_filter_q_reg_chain_5__2_), .A2(
        my_filter_delay_line_delay_chain_5_n48), .ZN(
        my_filter_delay_line_delay_chain_5_n82) );
  OAI21_X1 my_filter_delay_line_delay_chain_5_U11 ( .B1(
        my_filter_delay_line_delay_chain_5_n94), .B2(
        my_filter_delay_line_delay_chain_5_n77), .A(
        my_filter_delay_line_delay_chain_5_n82), .ZN(
        my_filter_delay_line_delay_chain_5_n54) );
  NAND2_X1 my_filter_delay_line_delay_chain_5_U10 ( .A1(
        my_filter_q_reg_chain_5__1_), .A2(
        my_filter_delay_line_delay_chain_5_n48), .ZN(
        my_filter_delay_line_delay_chain_5_n81) );
  OAI21_X1 my_filter_delay_line_delay_chain_5_U9 ( .B1(
        my_filter_delay_line_delay_chain_5_n94), .B2(
        my_filter_delay_line_delay_chain_5_n78), .A(
        my_filter_delay_line_delay_chain_5_n81), .ZN(
        my_filter_delay_line_delay_chain_5_n53) );
  NAND2_X1 my_filter_delay_line_delay_chain_5_U8 ( .A1(
        my_filter_q_reg_chain_5__0_), .A2(
        my_filter_delay_line_delay_chain_5_n48), .ZN(
        my_filter_delay_line_delay_chain_5_n80) );
  OAI21_X1 my_filter_delay_line_delay_chain_5_U7 ( .B1(
        my_filter_delay_line_delay_chain_5_n94), .B2(
        my_filter_delay_line_delay_chain_5_n79), .A(
        my_filter_delay_line_delay_chain_5_n80), .ZN(
        my_filter_delay_line_delay_chain_5_n52) );
  INV_X1 my_filter_delay_line_delay_chain_5_U6 ( .A(my_filter_delay_line_n8), 
        .ZN(my_filter_delay_line_delay_chain_5_n50) );
  INV_X1 my_filter_delay_line_delay_chain_5_U5 ( .A(
        my_filter_delay_line_delay_chain_5_n50), .ZN(
        my_filter_delay_line_delay_chain_5_n48) );
  NAND2_X1 my_filter_delay_line_delay_chain_5_U4 ( .A1(
        my_filter_delay_line_delay_chain_5_n51), .A2(
        my_filter_delay_line_delay_chain_5_n50), .ZN(
        my_filter_delay_line_delay_chain_5_n94) );
  BUF_X1 my_filter_delay_line_delay_chain_5_U3 ( .A(my_filter_delay_line_n13), 
        .Z(my_filter_delay_line_delay_chain_5_n51) );
  DFFR_X1 my_filter_delay_line_delay_chain_5_q_reg_0_ ( .D(
        my_filter_delay_line_delay_chain_5_n52), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_5_n51), .Q(
        my_filter_q_reg_chain_6__0_), .QN(
        my_filter_delay_line_delay_chain_5_n79) );
  DFFR_X1 my_filter_delay_line_delay_chain_5_q_reg_1_ ( .D(
        my_filter_delay_line_delay_chain_5_n53), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_5_n51), .Q(
        my_filter_q_reg_chain_6__1_), .QN(
        my_filter_delay_line_delay_chain_5_n78) );
  DFFR_X1 my_filter_delay_line_delay_chain_5_q_reg_2_ ( .D(
        my_filter_delay_line_delay_chain_5_n54), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_5_n51), .Q(
        my_filter_q_reg_chain_6__2_), .QN(
        my_filter_delay_line_delay_chain_5_n77) );
  DFFR_X1 my_filter_delay_line_delay_chain_5_q_reg_3_ ( .D(
        my_filter_delay_line_delay_chain_5_n55), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_5_n51), .Q(
        my_filter_q_reg_chain_6__3_), .QN(
        my_filter_delay_line_delay_chain_5_n76) );
  DFFR_X1 my_filter_delay_line_delay_chain_5_q_reg_4_ ( .D(
        my_filter_delay_line_delay_chain_5_n56), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_5_n51), .Q(
        my_filter_q_reg_chain_6__4_), .QN(
        my_filter_delay_line_delay_chain_5_n75) );
  DFFR_X1 my_filter_delay_line_delay_chain_5_q_reg_5_ ( .D(
        my_filter_delay_line_delay_chain_5_n57), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_5_n51), .Q(
        my_filter_q_reg_chain_6__5_), .QN(
        my_filter_delay_line_delay_chain_5_n74) );
  DFFR_X1 my_filter_delay_line_delay_chain_5_q_reg_6_ ( .D(
        my_filter_delay_line_delay_chain_5_n58), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_5_n51), .Q(
        my_filter_q_reg_chain_6__6_), .QN(
        my_filter_delay_line_delay_chain_5_n73) );
  DFFR_X1 my_filter_delay_line_delay_chain_5_q_reg_7_ ( .D(
        my_filter_delay_line_delay_chain_5_n59), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_5_n51), .Q(
        my_filter_q_reg_chain_6__7_), .QN(
        my_filter_delay_line_delay_chain_5_n72) );
  DFFR_X1 my_filter_delay_line_delay_chain_5_q_reg_8_ ( .D(
        my_filter_delay_line_delay_chain_5_n60), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_5_n51), .Q(
        my_filter_q_reg_chain_6__8_), .QN(
        my_filter_delay_line_delay_chain_5_n71) );
  DFFR_X1 my_filter_delay_line_delay_chain_5_q_reg_9_ ( .D(
        my_filter_delay_line_delay_chain_5_n61), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_5_n51), .Q(
        my_filter_q_reg_chain_6__9_), .QN(
        my_filter_delay_line_delay_chain_5_n70) );
  DFFR_X1 my_filter_delay_line_delay_chain_5_q_reg_10_ ( .D(
        my_filter_delay_line_delay_chain_5_n62), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_5_n51), .Q(
        my_filter_q_reg_chain_6__10_), .QN(
        my_filter_delay_line_delay_chain_5_n69) );
  DFFR_X1 my_filter_delay_line_delay_chain_5_q_reg_11_ ( .D(
        my_filter_delay_line_delay_chain_5_n63), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_5_n51), .Q(
        my_filter_q_reg_chain_6__11_), .QN(
        my_filter_delay_line_delay_chain_5_n68) );
  DFFR_X1 my_filter_delay_line_delay_chain_5_q_reg_12_ ( .D(
        my_filter_delay_line_delay_chain_5_n64), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_5_n51), .Q(
        my_filter_q_reg_chain_6__12_), .QN(
        my_filter_delay_line_delay_chain_5_n67) );
  DFFR_X1 my_filter_delay_line_delay_chain_5_q_reg_13_ ( .D(
        my_filter_delay_line_delay_chain_5_n65), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_5_n51), .Q(
        my_filter_q_reg_chain_6__13_), .QN(
        my_filter_delay_line_delay_chain_5_n66) );
  NAND2_X1 my_filter_delay_line_delay_chain_6_U34 ( .A1(
        my_filter_delay_line_n8), .A2(my_filter_q_reg_chain_6__13_), .ZN(
        my_filter_delay_line_delay_chain_6_n92) );
  OAI21_X1 my_filter_delay_line_delay_chain_6_U33 ( .B1(
        my_filter_delay_line_delay_chain_6_n93), .B2(
        my_filter_delay_line_delay_chain_6_n65), .A(
        my_filter_delay_line_delay_chain_6_n92), .ZN(
        my_filter_delay_line_delay_chain_6_n64) );
  NAND2_X1 my_filter_delay_line_delay_chain_6_U32 ( .A1(
        my_filter_q_reg_chain_6__12_), .A2(my_filter_delay_line_n8), .ZN(
        my_filter_delay_line_delay_chain_6_n91) );
  OAI21_X1 my_filter_delay_line_delay_chain_6_U31 ( .B1(
        my_filter_delay_line_delay_chain_6_n93), .B2(
        my_filter_delay_line_delay_chain_6_n66), .A(
        my_filter_delay_line_delay_chain_6_n91), .ZN(
        my_filter_delay_line_delay_chain_6_n63) );
  NAND2_X1 my_filter_delay_line_delay_chain_6_U30 ( .A1(
        my_filter_q_reg_chain_6__11_), .A2(
        my_filter_delay_line_delay_chain_6_n48), .ZN(
        my_filter_delay_line_delay_chain_6_n90) );
  OAI21_X1 my_filter_delay_line_delay_chain_6_U29 ( .B1(
        my_filter_delay_line_delay_chain_6_n93), .B2(
        my_filter_delay_line_delay_chain_6_n67), .A(
        my_filter_delay_line_delay_chain_6_n90), .ZN(
        my_filter_delay_line_delay_chain_6_n62) );
  NAND2_X1 my_filter_delay_line_delay_chain_6_U28 ( .A1(
        my_filter_q_reg_chain_6__10_), .A2(
        my_filter_delay_line_delay_chain_6_n48), .ZN(
        my_filter_delay_line_delay_chain_6_n89) );
  OAI21_X1 my_filter_delay_line_delay_chain_6_U27 ( .B1(
        my_filter_delay_line_delay_chain_6_n93), .B2(
        my_filter_delay_line_delay_chain_6_n68), .A(
        my_filter_delay_line_delay_chain_6_n89), .ZN(
        my_filter_delay_line_delay_chain_6_n61) );
  NAND2_X1 my_filter_delay_line_delay_chain_6_U26 ( .A1(
        my_filter_q_reg_chain_6__9_), .A2(
        my_filter_delay_line_delay_chain_6_n48), .ZN(
        my_filter_delay_line_delay_chain_6_n88) );
  OAI21_X1 my_filter_delay_line_delay_chain_6_U25 ( .B1(
        my_filter_delay_line_delay_chain_6_n93), .B2(
        my_filter_delay_line_delay_chain_6_n69), .A(
        my_filter_delay_line_delay_chain_6_n88), .ZN(
        my_filter_delay_line_delay_chain_6_n60) );
  NAND2_X1 my_filter_delay_line_delay_chain_6_U24 ( .A1(
        my_filter_q_reg_chain_6__8_), .A2(
        my_filter_delay_line_delay_chain_6_n48), .ZN(
        my_filter_delay_line_delay_chain_6_n87) );
  OAI21_X1 my_filter_delay_line_delay_chain_6_U23 ( .B1(
        my_filter_delay_line_delay_chain_6_n93), .B2(
        my_filter_delay_line_delay_chain_6_n70), .A(
        my_filter_delay_line_delay_chain_6_n87), .ZN(
        my_filter_delay_line_delay_chain_6_n59) );
  NAND2_X1 my_filter_delay_line_delay_chain_6_U22 ( .A1(
        my_filter_q_reg_chain_6__7_), .A2(
        my_filter_delay_line_delay_chain_6_n48), .ZN(
        my_filter_delay_line_delay_chain_6_n86) );
  OAI21_X1 my_filter_delay_line_delay_chain_6_U21 ( .B1(
        my_filter_delay_line_delay_chain_6_n93), .B2(
        my_filter_delay_line_delay_chain_6_n71), .A(
        my_filter_delay_line_delay_chain_6_n86), .ZN(
        my_filter_delay_line_delay_chain_6_n58) );
  NAND2_X1 my_filter_delay_line_delay_chain_6_U20 ( .A1(
        my_filter_q_reg_chain_6__6_), .A2(
        my_filter_delay_line_delay_chain_6_n48), .ZN(
        my_filter_delay_line_delay_chain_6_n85) );
  OAI21_X1 my_filter_delay_line_delay_chain_6_U19 ( .B1(
        my_filter_delay_line_delay_chain_6_n93), .B2(
        my_filter_delay_line_delay_chain_6_n72), .A(
        my_filter_delay_line_delay_chain_6_n85), .ZN(
        my_filter_delay_line_delay_chain_6_n57) );
  NAND2_X1 my_filter_delay_line_delay_chain_6_U18 ( .A1(
        my_filter_q_reg_chain_6__5_), .A2(
        my_filter_delay_line_delay_chain_6_n48), .ZN(
        my_filter_delay_line_delay_chain_6_n84) );
  OAI21_X1 my_filter_delay_line_delay_chain_6_U17 ( .B1(
        my_filter_delay_line_delay_chain_6_n93), .B2(
        my_filter_delay_line_delay_chain_6_n73), .A(
        my_filter_delay_line_delay_chain_6_n84), .ZN(
        my_filter_delay_line_delay_chain_6_n56) );
  NAND2_X1 my_filter_delay_line_delay_chain_6_U16 ( .A1(
        my_filter_q_reg_chain_6__4_), .A2(
        my_filter_delay_line_delay_chain_6_n48), .ZN(
        my_filter_delay_line_delay_chain_6_n83) );
  OAI21_X1 my_filter_delay_line_delay_chain_6_U15 ( .B1(
        my_filter_delay_line_delay_chain_6_n93), .B2(
        my_filter_delay_line_delay_chain_6_n74), .A(
        my_filter_delay_line_delay_chain_6_n83), .ZN(
        my_filter_delay_line_delay_chain_6_n55) );
  NAND2_X1 my_filter_delay_line_delay_chain_6_U14 ( .A1(
        my_filter_q_reg_chain_6__3_), .A2(
        my_filter_delay_line_delay_chain_6_n48), .ZN(
        my_filter_delay_line_delay_chain_6_n82) );
  OAI21_X1 my_filter_delay_line_delay_chain_6_U13 ( .B1(
        my_filter_delay_line_delay_chain_6_n93), .B2(
        my_filter_delay_line_delay_chain_6_n75), .A(
        my_filter_delay_line_delay_chain_6_n82), .ZN(
        my_filter_delay_line_delay_chain_6_n54) );
  NAND2_X1 my_filter_delay_line_delay_chain_6_U12 ( .A1(
        my_filter_q_reg_chain_6__2_), .A2(
        my_filter_delay_line_delay_chain_6_n48), .ZN(
        my_filter_delay_line_delay_chain_6_n81) );
  OAI21_X1 my_filter_delay_line_delay_chain_6_U11 ( .B1(
        my_filter_delay_line_delay_chain_6_n93), .B2(
        my_filter_delay_line_delay_chain_6_n76), .A(
        my_filter_delay_line_delay_chain_6_n81), .ZN(
        my_filter_delay_line_delay_chain_6_n53) );
  NAND2_X1 my_filter_delay_line_delay_chain_6_U10 ( .A1(
        my_filter_q_reg_chain_6__1_), .A2(
        my_filter_delay_line_delay_chain_6_n48), .ZN(
        my_filter_delay_line_delay_chain_6_n80) );
  OAI21_X1 my_filter_delay_line_delay_chain_6_U9 ( .B1(
        my_filter_delay_line_delay_chain_6_n93), .B2(
        my_filter_delay_line_delay_chain_6_n77), .A(
        my_filter_delay_line_delay_chain_6_n80), .ZN(
        my_filter_delay_line_delay_chain_6_n52) );
  NAND2_X1 my_filter_delay_line_delay_chain_6_U8 ( .A1(
        my_filter_q_reg_chain_6__0_), .A2(
        my_filter_delay_line_delay_chain_6_n48), .ZN(
        my_filter_delay_line_delay_chain_6_n79) );
  OAI21_X1 my_filter_delay_line_delay_chain_6_U7 ( .B1(
        my_filter_delay_line_delay_chain_6_n93), .B2(
        my_filter_delay_line_delay_chain_6_n78), .A(
        my_filter_delay_line_delay_chain_6_n79), .ZN(
        my_filter_delay_line_delay_chain_6_n51) );
  INV_X1 my_filter_delay_line_delay_chain_6_U6 ( .A(my_filter_delay_line_n8), 
        .ZN(my_filter_delay_line_delay_chain_6_n49) );
  INV_X1 my_filter_delay_line_delay_chain_6_U5 ( .A(
        my_filter_delay_line_delay_chain_6_n49), .ZN(
        my_filter_delay_line_delay_chain_6_n48) );
  NAND2_X1 my_filter_delay_line_delay_chain_6_U4 ( .A1(
        my_filter_delay_line_delay_chain_6_n50), .A2(
        my_filter_delay_line_delay_chain_6_n49), .ZN(
        my_filter_delay_line_delay_chain_6_n93) );
  BUF_X1 my_filter_delay_line_delay_chain_6_U3 ( .A(my_filter_delay_line_n13), 
        .Z(my_filter_delay_line_delay_chain_6_n50) );
  DFFR_X1 my_filter_delay_line_delay_chain_6_q_reg_0_ ( .D(
        my_filter_delay_line_delay_chain_6_n51), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_6_n50), .Q(
        my_filter_q_reg_chain_7__0_), .QN(
        my_filter_delay_line_delay_chain_6_n78) );
  DFFR_X1 my_filter_delay_line_delay_chain_6_q_reg_1_ ( .D(
        my_filter_delay_line_delay_chain_6_n52), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_6_n50), .Q(
        my_filter_q_reg_chain_7__1_), .QN(
        my_filter_delay_line_delay_chain_6_n77) );
  DFFR_X1 my_filter_delay_line_delay_chain_6_q_reg_2_ ( .D(
        my_filter_delay_line_delay_chain_6_n53), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_6_n50), .Q(
        my_filter_q_reg_chain_7__2_), .QN(
        my_filter_delay_line_delay_chain_6_n76) );
  DFFR_X1 my_filter_delay_line_delay_chain_6_q_reg_3_ ( .D(
        my_filter_delay_line_delay_chain_6_n54), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_6_n50), .Q(
        my_filter_q_reg_chain_7__3_), .QN(
        my_filter_delay_line_delay_chain_6_n75) );
  DFFR_X1 my_filter_delay_line_delay_chain_6_q_reg_4_ ( .D(
        my_filter_delay_line_delay_chain_6_n55), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_6_n50), .Q(
        my_filter_q_reg_chain_7__4_), .QN(
        my_filter_delay_line_delay_chain_6_n74) );
  DFFR_X1 my_filter_delay_line_delay_chain_6_q_reg_5_ ( .D(
        my_filter_delay_line_delay_chain_6_n56), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_6_n50), .Q(
        my_filter_q_reg_chain_7__5_), .QN(
        my_filter_delay_line_delay_chain_6_n73) );
  DFFR_X1 my_filter_delay_line_delay_chain_6_q_reg_6_ ( .D(
        my_filter_delay_line_delay_chain_6_n57), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_6_n50), .Q(
        my_filter_q_reg_chain_7__6_), .QN(
        my_filter_delay_line_delay_chain_6_n72) );
  DFFR_X1 my_filter_delay_line_delay_chain_6_q_reg_7_ ( .D(
        my_filter_delay_line_delay_chain_6_n58), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_6_n50), .Q(
        my_filter_q_reg_chain_7__7_), .QN(
        my_filter_delay_line_delay_chain_6_n71) );
  DFFR_X1 my_filter_delay_line_delay_chain_6_q_reg_8_ ( .D(
        my_filter_delay_line_delay_chain_6_n59), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_6_n50), .Q(
        my_filter_q_reg_chain_7__8_), .QN(
        my_filter_delay_line_delay_chain_6_n70) );
  DFFR_X1 my_filter_delay_line_delay_chain_6_q_reg_9_ ( .D(
        my_filter_delay_line_delay_chain_6_n60), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_6_n50), .Q(
        my_filter_q_reg_chain_7__9_), .QN(
        my_filter_delay_line_delay_chain_6_n69) );
  DFFR_X1 my_filter_delay_line_delay_chain_6_q_reg_10_ ( .D(
        my_filter_delay_line_delay_chain_6_n61), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_6_n50), .Q(
        my_filter_q_reg_chain_7__10_), .QN(
        my_filter_delay_line_delay_chain_6_n68) );
  DFFR_X1 my_filter_delay_line_delay_chain_6_q_reg_11_ ( .D(
        my_filter_delay_line_delay_chain_6_n62), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_6_n50), .Q(
        my_filter_q_reg_chain_7__11_), .QN(
        my_filter_delay_line_delay_chain_6_n67) );
  DFFR_X1 my_filter_delay_line_delay_chain_6_q_reg_12_ ( .D(
        my_filter_delay_line_delay_chain_6_n63), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_6_n50), .Q(
        my_filter_q_reg_chain_7__12_), .QN(
        my_filter_delay_line_delay_chain_6_n66) );
  DFFR_X1 my_filter_delay_line_delay_chain_6_q_reg_13_ ( .D(
        my_filter_delay_line_delay_chain_6_n64), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_6_n50), .Q(
        my_filter_q_reg_chain_7__13_), .QN(
        my_filter_delay_line_delay_chain_6_n65) );
  NAND2_X1 my_filter_delay_line_delay_chain_7_U34 ( .A1(
        my_filter_delay_line_n8), .A2(my_filter_q_reg_chain_7__13_), .ZN(
        my_filter_delay_line_delay_chain_7_n92) );
  OAI21_X1 my_filter_delay_line_delay_chain_7_U33 ( .B1(
        my_filter_delay_line_delay_chain_7_n93), .B2(
        my_filter_delay_line_delay_chain_7_n65), .A(
        my_filter_delay_line_delay_chain_7_n92), .ZN(
        my_filter_delay_line_delay_chain_7_n64) );
  NAND2_X1 my_filter_delay_line_delay_chain_7_U32 ( .A1(
        my_filter_q_reg_chain_7__12_), .A2(my_filter_delay_line_n8), .ZN(
        my_filter_delay_line_delay_chain_7_n91) );
  OAI21_X1 my_filter_delay_line_delay_chain_7_U31 ( .B1(
        my_filter_delay_line_delay_chain_7_n93), .B2(
        my_filter_delay_line_delay_chain_7_n66), .A(
        my_filter_delay_line_delay_chain_7_n91), .ZN(
        my_filter_delay_line_delay_chain_7_n63) );
  NAND2_X1 my_filter_delay_line_delay_chain_7_U30 ( .A1(
        my_filter_q_reg_chain_7__11_), .A2(
        my_filter_delay_line_delay_chain_7_n48), .ZN(
        my_filter_delay_line_delay_chain_7_n90) );
  OAI21_X1 my_filter_delay_line_delay_chain_7_U29 ( .B1(
        my_filter_delay_line_delay_chain_7_n93), .B2(
        my_filter_delay_line_delay_chain_7_n67), .A(
        my_filter_delay_line_delay_chain_7_n90), .ZN(
        my_filter_delay_line_delay_chain_7_n62) );
  NAND2_X1 my_filter_delay_line_delay_chain_7_U28 ( .A1(
        my_filter_q_reg_chain_7__10_), .A2(
        my_filter_delay_line_delay_chain_7_n48), .ZN(
        my_filter_delay_line_delay_chain_7_n89) );
  OAI21_X1 my_filter_delay_line_delay_chain_7_U27 ( .B1(
        my_filter_delay_line_delay_chain_7_n93), .B2(
        my_filter_delay_line_delay_chain_7_n68), .A(
        my_filter_delay_line_delay_chain_7_n89), .ZN(
        my_filter_delay_line_delay_chain_7_n61) );
  NAND2_X1 my_filter_delay_line_delay_chain_7_U26 ( .A1(
        my_filter_q_reg_chain_7__9_), .A2(
        my_filter_delay_line_delay_chain_7_n48), .ZN(
        my_filter_delay_line_delay_chain_7_n88) );
  OAI21_X1 my_filter_delay_line_delay_chain_7_U25 ( .B1(
        my_filter_delay_line_delay_chain_7_n93), .B2(
        my_filter_delay_line_delay_chain_7_n69), .A(
        my_filter_delay_line_delay_chain_7_n88), .ZN(
        my_filter_delay_line_delay_chain_7_n60) );
  NAND2_X1 my_filter_delay_line_delay_chain_7_U24 ( .A1(
        my_filter_q_reg_chain_7__8_), .A2(
        my_filter_delay_line_delay_chain_7_n48), .ZN(
        my_filter_delay_line_delay_chain_7_n87) );
  OAI21_X1 my_filter_delay_line_delay_chain_7_U23 ( .B1(
        my_filter_delay_line_delay_chain_7_n93), .B2(
        my_filter_delay_line_delay_chain_7_n70), .A(
        my_filter_delay_line_delay_chain_7_n87), .ZN(
        my_filter_delay_line_delay_chain_7_n59) );
  NAND2_X1 my_filter_delay_line_delay_chain_7_U22 ( .A1(
        my_filter_q_reg_chain_7__7_), .A2(
        my_filter_delay_line_delay_chain_7_n48), .ZN(
        my_filter_delay_line_delay_chain_7_n86) );
  OAI21_X1 my_filter_delay_line_delay_chain_7_U21 ( .B1(
        my_filter_delay_line_delay_chain_7_n93), .B2(
        my_filter_delay_line_delay_chain_7_n71), .A(
        my_filter_delay_line_delay_chain_7_n86), .ZN(
        my_filter_delay_line_delay_chain_7_n58) );
  NAND2_X1 my_filter_delay_line_delay_chain_7_U20 ( .A1(
        my_filter_q_reg_chain_7__6_), .A2(
        my_filter_delay_line_delay_chain_7_n48), .ZN(
        my_filter_delay_line_delay_chain_7_n85) );
  OAI21_X1 my_filter_delay_line_delay_chain_7_U19 ( .B1(
        my_filter_delay_line_delay_chain_7_n93), .B2(
        my_filter_delay_line_delay_chain_7_n72), .A(
        my_filter_delay_line_delay_chain_7_n85), .ZN(
        my_filter_delay_line_delay_chain_7_n57) );
  NAND2_X1 my_filter_delay_line_delay_chain_7_U18 ( .A1(
        my_filter_q_reg_chain_7__5_), .A2(
        my_filter_delay_line_delay_chain_7_n48), .ZN(
        my_filter_delay_line_delay_chain_7_n84) );
  OAI21_X1 my_filter_delay_line_delay_chain_7_U17 ( .B1(
        my_filter_delay_line_delay_chain_7_n93), .B2(
        my_filter_delay_line_delay_chain_7_n73), .A(
        my_filter_delay_line_delay_chain_7_n84), .ZN(
        my_filter_delay_line_delay_chain_7_n56) );
  NAND2_X1 my_filter_delay_line_delay_chain_7_U16 ( .A1(
        my_filter_q_reg_chain_7__4_), .A2(
        my_filter_delay_line_delay_chain_7_n48), .ZN(
        my_filter_delay_line_delay_chain_7_n83) );
  OAI21_X1 my_filter_delay_line_delay_chain_7_U15 ( .B1(
        my_filter_delay_line_delay_chain_7_n93), .B2(
        my_filter_delay_line_delay_chain_7_n74), .A(
        my_filter_delay_line_delay_chain_7_n83), .ZN(
        my_filter_delay_line_delay_chain_7_n55) );
  NAND2_X1 my_filter_delay_line_delay_chain_7_U14 ( .A1(
        my_filter_q_reg_chain_7__3_), .A2(
        my_filter_delay_line_delay_chain_7_n48), .ZN(
        my_filter_delay_line_delay_chain_7_n82) );
  OAI21_X1 my_filter_delay_line_delay_chain_7_U13 ( .B1(
        my_filter_delay_line_delay_chain_7_n93), .B2(
        my_filter_delay_line_delay_chain_7_n75), .A(
        my_filter_delay_line_delay_chain_7_n82), .ZN(
        my_filter_delay_line_delay_chain_7_n54) );
  NAND2_X1 my_filter_delay_line_delay_chain_7_U12 ( .A1(
        my_filter_q_reg_chain_7__2_), .A2(
        my_filter_delay_line_delay_chain_7_n48), .ZN(
        my_filter_delay_line_delay_chain_7_n81) );
  OAI21_X1 my_filter_delay_line_delay_chain_7_U11 ( .B1(
        my_filter_delay_line_delay_chain_7_n93), .B2(
        my_filter_delay_line_delay_chain_7_n76), .A(
        my_filter_delay_line_delay_chain_7_n81), .ZN(
        my_filter_delay_line_delay_chain_7_n53) );
  NAND2_X1 my_filter_delay_line_delay_chain_7_U10 ( .A1(
        my_filter_q_reg_chain_7__1_), .A2(
        my_filter_delay_line_delay_chain_7_n48), .ZN(
        my_filter_delay_line_delay_chain_7_n80) );
  OAI21_X1 my_filter_delay_line_delay_chain_7_U9 ( .B1(
        my_filter_delay_line_delay_chain_7_n93), .B2(
        my_filter_delay_line_delay_chain_7_n77), .A(
        my_filter_delay_line_delay_chain_7_n80), .ZN(
        my_filter_delay_line_delay_chain_7_n52) );
  NAND2_X1 my_filter_delay_line_delay_chain_7_U8 ( .A1(
        my_filter_q_reg_chain_7__0_), .A2(
        my_filter_delay_line_delay_chain_7_n48), .ZN(
        my_filter_delay_line_delay_chain_7_n79) );
  OAI21_X1 my_filter_delay_line_delay_chain_7_U7 ( .B1(
        my_filter_delay_line_delay_chain_7_n93), .B2(
        my_filter_delay_line_delay_chain_7_n78), .A(
        my_filter_delay_line_delay_chain_7_n79), .ZN(
        my_filter_delay_line_delay_chain_7_n51) );
  INV_X1 my_filter_delay_line_delay_chain_7_U6 ( .A(my_filter_delay_line_n8), 
        .ZN(my_filter_delay_line_delay_chain_7_n49) );
  INV_X1 my_filter_delay_line_delay_chain_7_U5 ( .A(
        my_filter_delay_line_delay_chain_7_n49), .ZN(
        my_filter_delay_line_delay_chain_7_n48) );
  NAND2_X1 my_filter_delay_line_delay_chain_7_U4 ( .A1(
        my_filter_delay_line_delay_chain_7_n50), .A2(
        my_filter_delay_line_delay_chain_7_n49), .ZN(
        my_filter_delay_line_delay_chain_7_n93) );
  BUF_X1 my_filter_delay_line_delay_chain_7_U3 ( .A(my_filter_delay_line_n14), 
        .Z(my_filter_delay_line_delay_chain_7_n50) );
  DFFR_X1 my_filter_delay_line_delay_chain_7_q_reg_0_ ( .D(
        my_filter_delay_line_delay_chain_7_n51), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_7_n50), .Q(
        my_filter_q_reg_chain_8__0_), .QN(
        my_filter_delay_line_delay_chain_7_n78) );
  DFFR_X1 my_filter_delay_line_delay_chain_7_q_reg_1_ ( .D(
        my_filter_delay_line_delay_chain_7_n52), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_7_n50), .Q(
        my_filter_q_reg_chain_8__1_), .QN(
        my_filter_delay_line_delay_chain_7_n77) );
  DFFR_X1 my_filter_delay_line_delay_chain_7_q_reg_2_ ( .D(
        my_filter_delay_line_delay_chain_7_n53), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_7_n50), .Q(
        my_filter_q_reg_chain_8__2_), .QN(
        my_filter_delay_line_delay_chain_7_n76) );
  DFFR_X1 my_filter_delay_line_delay_chain_7_q_reg_3_ ( .D(
        my_filter_delay_line_delay_chain_7_n54), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_7_n50), .Q(
        my_filter_q_reg_chain_8__3_), .QN(
        my_filter_delay_line_delay_chain_7_n75) );
  DFFR_X1 my_filter_delay_line_delay_chain_7_q_reg_4_ ( .D(
        my_filter_delay_line_delay_chain_7_n55), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_7_n50), .Q(
        my_filter_q_reg_chain_8__4_), .QN(
        my_filter_delay_line_delay_chain_7_n74) );
  DFFR_X1 my_filter_delay_line_delay_chain_7_q_reg_5_ ( .D(
        my_filter_delay_line_delay_chain_7_n56), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_7_n50), .Q(
        my_filter_q_reg_chain_8__5_), .QN(
        my_filter_delay_line_delay_chain_7_n73) );
  DFFR_X1 my_filter_delay_line_delay_chain_7_q_reg_6_ ( .D(
        my_filter_delay_line_delay_chain_7_n57), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_7_n50), .Q(
        my_filter_q_reg_chain_8__6_), .QN(
        my_filter_delay_line_delay_chain_7_n72) );
  DFFR_X1 my_filter_delay_line_delay_chain_7_q_reg_7_ ( .D(
        my_filter_delay_line_delay_chain_7_n58), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_7_n50), .Q(
        my_filter_q_reg_chain_8__7_), .QN(
        my_filter_delay_line_delay_chain_7_n71) );
  DFFR_X1 my_filter_delay_line_delay_chain_7_q_reg_8_ ( .D(
        my_filter_delay_line_delay_chain_7_n59), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_7_n50), .Q(
        my_filter_q_reg_chain_8__8_), .QN(
        my_filter_delay_line_delay_chain_7_n70) );
  DFFR_X1 my_filter_delay_line_delay_chain_7_q_reg_9_ ( .D(
        my_filter_delay_line_delay_chain_7_n60), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_7_n50), .Q(
        my_filter_q_reg_chain_8__9_), .QN(
        my_filter_delay_line_delay_chain_7_n69) );
  DFFR_X1 my_filter_delay_line_delay_chain_7_q_reg_10_ ( .D(
        my_filter_delay_line_delay_chain_7_n61), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_7_n50), .Q(
        my_filter_q_reg_chain_8__10_), .QN(
        my_filter_delay_line_delay_chain_7_n68) );
  DFFR_X1 my_filter_delay_line_delay_chain_7_q_reg_11_ ( .D(
        my_filter_delay_line_delay_chain_7_n62), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_7_n50), .Q(
        my_filter_q_reg_chain_8__11_), .QN(
        my_filter_delay_line_delay_chain_7_n67) );
  DFFR_X1 my_filter_delay_line_delay_chain_7_q_reg_12_ ( .D(
        my_filter_delay_line_delay_chain_7_n63), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_7_n50), .Q(
        my_filter_q_reg_chain_8__12_), .QN(
        my_filter_delay_line_delay_chain_7_n66) );
  DFFR_X1 my_filter_delay_line_delay_chain_7_q_reg_13_ ( .D(
        my_filter_delay_line_delay_chain_7_n64), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_7_n50), .Q(
        my_filter_q_reg_chain_8__13_), .QN(
        my_filter_delay_line_delay_chain_7_n65) );
  NAND2_X1 my_filter_delay_line_delay_chain_8_U34 ( .A1(
        my_filter_delay_line_n8), .A2(my_filter_q_reg_chain_8__13_), .ZN(
        my_filter_delay_line_delay_chain_8_n92) );
  OAI21_X1 my_filter_delay_line_delay_chain_8_U33 ( .B1(
        my_filter_delay_line_delay_chain_8_n93), .B2(
        my_filter_delay_line_delay_chain_8_n65), .A(
        my_filter_delay_line_delay_chain_8_n92), .ZN(
        my_filter_delay_line_delay_chain_8_n64) );
  NAND2_X1 my_filter_delay_line_delay_chain_8_U32 ( .A1(
        my_filter_q_reg_chain_8__12_), .A2(my_filter_delay_line_n8), .ZN(
        my_filter_delay_line_delay_chain_8_n91) );
  OAI21_X1 my_filter_delay_line_delay_chain_8_U31 ( .B1(
        my_filter_delay_line_delay_chain_8_n93), .B2(
        my_filter_delay_line_delay_chain_8_n66), .A(
        my_filter_delay_line_delay_chain_8_n91), .ZN(
        my_filter_delay_line_delay_chain_8_n63) );
  NAND2_X1 my_filter_delay_line_delay_chain_8_U30 ( .A1(
        my_filter_q_reg_chain_8__11_), .A2(
        my_filter_delay_line_delay_chain_8_n48), .ZN(
        my_filter_delay_line_delay_chain_8_n90) );
  OAI21_X1 my_filter_delay_line_delay_chain_8_U29 ( .B1(
        my_filter_delay_line_delay_chain_8_n93), .B2(
        my_filter_delay_line_delay_chain_8_n67), .A(
        my_filter_delay_line_delay_chain_8_n90), .ZN(
        my_filter_delay_line_delay_chain_8_n62) );
  NAND2_X1 my_filter_delay_line_delay_chain_8_U28 ( .A1(
        my_filter_q_reg_chain_8__10_), .A2(
        my_filter_delay_line_delay_chain_8_n48), .ZN(
        my_filter_delay_line_delay_chain_8_n89) );
  OAI21_X1 my_filter_delay_line_delay_chain_8_U27 ( .B1(
        my_filter_delay_line_delay_chain_8_n93), .B2(
        my_filter_delay_line_delay_chain_8_n68), .A(
        my_filter_delay_line_delay_chain_8_n89), .ZN(
        my_filter_delay_line_delay_chain_8_n61) );
  NAND2_X1 my_filter_delay_line_delay_chain_8_U26 ( .A1(
        my_filter_q_reg_chain_8__9_), .A2(
        my_filter_delay_line_delay_chain_8_n48), .ZN(
        my_filter_delay_line_delay_chain_8_n88) );
  OAI21_X1 my_filter_delay_line_delay_chain_8_U25 ( .B1(
        my_filter_delay_line_delay_chain_8_n93), .B2(
        my_filter_delay_line_delay_chain_8_n69), .A(
        my_filter_delay_line_delay_chain_8_n88), .ZN(
        my_filter_delay_line_delay_chain_8_n60) );
  NAND2_X1 my_filter_delay_line_delay_chain_8_U24 ( .A1(
        my_filter_q_reg_chain_8__8_), .A2(
        my_filter_delay_line_delay_chain_8_n48), .ZN(
        my_filter_delay_line_delay_chain_8_n87) );
  OAI21_X1 my_filter_delay_line_delay_chain_8_U23 ( .B1(
        my_filter_delay_line_delay_chain_8_n93), .B2(
        my_filter_delay_line_delay_chain_8_n70), .A(
        my_filter_delay_line_delay_chain_8_n87), .ZN(
        my_filter_delay_line_delay_chain_8_n59) );
  NAND2_X1 my_filter_delay_line_delay_chain_8_U22 ( .A1(
        my_filter_q_reg_chain_8__7_), .A2(
        my_filter_delay_line_delay_chain_8_n48), .ZN(
        my_filter_delay_line_delay_chain_8_n86) );
  OAI21_X1 my_filter_delay_line_delay_chain_8_U21 ( .B1(
        my_filter_delay_line_delay_chain_8_n93), .B2(
        my_filter_delay_line_delay_chain_8_n71), .A(
        my_filter_delay_line_delay_chain_8_n86), .ZN(
        my_filter_delay_line_delay_chain_8_n58) );
  NAND2_X1 my_filter_delay_line_delay_chain_8_U20 ( .A1(
        my_filter_q_reg_chain_8__6_), .A2(
        my_filter_delay_line_delay_chain_8_n48), .ZN(
        my_filter_delay_line_delay_chain_8_n85) );
  OAI21_X1 my_filter_delay_line_delay_chain_8_U19 ( .B1(
        my_filter_delay_line_delay_chain_8_n93), .B2(
        my_filter_delay_line_delay_chain_8_n72), .A(
        my_filter_delay_line_delay_chain_8_n85), .ZN(
        my_filter_delay_line_delay_chain_8_n57) );
  NAND2_X1 my_filter_delay_line_delay_chain_8_U18 ( .A1(
        my_filter_q_reg_chain_8__5_), .A2(
        my_filter_delay_line_delay_chain_8_n48), .ZN(
        my_filter_delay_line_delay_chain_8_n84) );
  OAI21_X1 my_filter_delay_line_delay_chain_8_U17 ( .B1(
        my_filter_delay_line_delay_chain_8_n93), .B2(
        my_filter_delay_line_delay_chain_8_n73), .A(
        my_filter_delay_line_delay_chain_8_n84), .ZN(
        my_filter_delay_line_delay_chain_8_n56) );
  NAND2_X1 my_filter_delay_line_delay_chain_8_U16 ( .A1(
        my_filter_q_reg_chain_8__4_), .A2(
        my_filter_delay_line_delay_chain_8_n48), .ZN(
        my_filter_delay_line_delay_chain_8_n83) );
  OAI21_X1 my_filter_delay_line_delay_chain_8_U15 ( .B1(
        my_filter_delay_line_delay_chain_8_n93), .B2(
        my_filter_delay_line_delay_chain_8_n74), .A(
        my_filter_delay_line_delay_chain_8_n83), .ZN(
        my_filter_delay_line_delay_chain_8_n55) );
  NAND2_X1 my_filter_delay_line_delay_chain_8_U14 ( .A1(
        my_filter_q_reg_chain_8__3_), .A2(
        my_filter_delay_line_delay_chain_8_n48), .ZN(
        my_filter_delay_line_delay_chain_8_n82) );
  OAI21_X1 my_filter_delay_line_delay_chain_8_U13 ( .B1(
        my_filter_delay_line_delay_chain_8_n93), .B2(
        my_filter_delay_line_delay_chain_8_n75), .A(
        my_filter_delay_line_delay_chain_8_n82), .ZN(
        my_filter_delay_line_delay_chain_8_n54) );
  NAND2_X1 my_filter_delay_line_delay_chain_8_U12 ( .A1(
        my_filter_q_reg_chain_8__2_), .A2(
        my_filter_delay_line_delay_chain_8_n48), .ZN(
        my_filter_delay_line_delay_chain_8_n81) );
  OAI21_X1 my_filter_delay_line_delay_chain_8_U11 ( .B1(
        my_filter_delay_line_delay_chain_8_n93), .B2(
        my_filter_delay_line_delay_chain_8_n76), .A(
        my_filter_delay_line_delay_chain_8_n81), .ZN(
        my_filter_delay_line_delay_chain_8_n53) );
  NAND2_X1 my_filter_delay_line_delay_chain_8_U10 ( .A1(
        my_filter_q_reg_chain_8__1_), .A2(
        my_filter_delay_line_delay_chain_8_n48), .ZN(
        my_filter_delay_line_delay_chain_8_n80) );
  OAI21_X1 my_filter_delay_line_delay_chain_8_U9 ( .B1(
        my_filter_delay_line_delay_chain_8_n93), .B2(
        my_filter_delay_line_delay_chain_8_n77), .A(
        my_filter_delay_line_delay_chain_8_n80), .ZN(
        my_filter_delay_line_delay_chain_8_n52) );
  NAND2_X1 my_filter_delay_line_delay_chain_8_U8 ( .A1(
        my_filter_q_reg_chain_8__0_), .A2(
        my_filter_delay_line_delay_chain_8_n48), .ZN(
        my_filter_delay_line_delay_chain_8_n79) );
  OAI21_X1 my_filter_delay_line_delay_chain_8_U7 ( .B1(
        my_filter_delay_line_delay_chain_8_n93), .B2(
        my_filter_delay_line_delay_chain_8_n78), .A(
        my_filter_delay_line_delay_chain_8_n79), .ZN(
        my_filter_delay_line_delay_chain_8_n51) );
  INV_X1 my_filter_delay_line_delay_chain_8_U6 ( .A(my_filter_delay_line_n8), 
        .ZN(my_filter_delay_line_delay_chain_8_n49) );
  INV_X1 my_filter_delay_line_delay_chain_8_U5 ( .A(
        my_filter_delay_line_delay_chain_8_n49), .ZN(
        my_filter_delay_line_delay_chain_8_n48) );
  NAND2_X1 my_filter_delay_line_delay_chain_8_U4 ( .A1(
        my_filter_delay_line_delay_chain_8_n50), .A2(
        my_filter_delay_line_delay_chain_8_n49), .ZN(
        my_filter_delay_line_delay_chain_8_n93) );
  BUF_X1 my_filter_delay_line_delay_chain_8_U3 ( .A(my_filter_delay_line_n14), 
        .Z(my_filter_delay_line_delay_chain_8_n50) );
  DFFR_X1 my_filter_delay_line_delay_chain_8_q_reg_0_ ( .D(
        my_filter_delay_line_delay_chain_8_n51), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_8_n50), .Q(
        my_filter_q_reg_chain_9__0_), .QN(
        my_filter_delay_line_delay_chain_8_n78) );
  DFFR_X1 my_filter_delay_line_delay_chain_8_q_reg_1_ ( .D(
        my_filter_delay_line_delay_chain_8_n52), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_8_n50), .Q(
        my_filter_q_reg_chain_9__1_), .QN(
        my_filter_delay_line_delay_chain_8_n77) );
  DFFR_X1 my_filter_delay_line_delay_chain_8_q_reg_2_ ( .D(
        my_filter_delay_line_delay_chain_8_n53), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_8_n50), .Q(
        my_filter_q_reg_chain_9__2_), .QN(
        my_filter_delay_line_delay_chain_8_n76) );
  DFFR_X1 my_filter_delay_line_delay_chain_8_q_reg_3_ ( .D(
        my_filter_delay_line_delay_chain_8_n54), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_8_n50), .Q(
        my_filter_q_reg_chain_9__3_), .QN(
        my_filter_delay_line_delay_chain_8_n75) );
  DFFR_X1 my_filter_delay_line_delay_chain_8_q_reg_4_ ( .D(
        my_filter_delay_line_delay_chain_8_n55), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_8_n50), .Q(
        my_filter_q_reg_chain_9__4_), .QN(
        my_filter_delay_line_delay_chain_8_n74) );
  DFFR_X1 my_filter_delay_line_delay_chain_8_q_reg_5_ ( .D(
        my_filter_delay_line_delay_chain_8_n56), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_8_n50), .Q(
        my_filter_q_reg_chain_9__5_), .QN(
        my_filter_delay_line_delay_chain_8_n73) );
  DFFR_X1 my_filter_delay_line_delay_chain_8_q_reg_6_ ( .D(
        my_filter_delay_line_delay_chain_8_n57), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_8_n50), .Q(
        my_filter_q_reg_chain_9__6_), .QN(
        my_filter_delay_line_delay_chain_8_n72) );
  DFFR_X1 my_filter_delay_line_delay_chain_8_q_reg_7_ ( .D(
        my_filter_delay_line_delay_chain_8_n58), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_8_n50), .Q(
        my_filter_q_reg_chain_9__7_), .QN(
        my_filter_delay_line_delay_chain_8_n71) );
  DFFR_X1 my_filter_delay_line_delay_chain_8_q_reg_8_ ( .D(
        my_filter_delay_line_delay_chain_8_n59), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_8_n50), .Q(
        my_filter_q_reg_chain_9__8_), .QN(
        my_filter_delay_line_delay_chain_8_n70) );
  DFFR_X1 my_filter_delay_line_delay_chain_8_q_reg_9_ ( .D(
        my_filter_delay_line_delay_chain_8_n60), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_8_n50), .Q(
        my_filter_q_reg_chain_9__9_), .QN(
        my_filter_delay_line_delay_chain_8_n69) );
  DFFR_X1 my_filter_delay_line_delay_chain_8_q_reg_10_ ( .D(
        my_filter_delay_line_delay_chain_8_n61), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_8_n50), .Q(
        my_filter_q_reg_chain_9__10_), .QN(
        my_filter_delay_line_delay_chain_8_n68) );
  DFFR_X1 my_filter_delay_line_delay_chain_8_q_reg_11_ ( .D(
        my_filter_delay_line_delay_chain_8_n62), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_8_n50), .Q(
        my_filter_q_reg_chain_9__11_), .QN(
        my_filter_delay_line_delay_chain_8_n67) );
  DFFR_X1 my_filter_delay_line_delay_chain_8_q_reg_12_ ( .D(
        my_filter_delay_line_delay_chain_8_n63), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_8_n50), .Q(
        my_filter_q_reg_chain_9__12_), .QN(
        my_filter_delay_line_delay_chain_8_n66) );
  DFFR_X1 my_filter_delay_line_delay_chain_8_q_reg_13_ ( .D(
        my_filter_delay_line_delay_chain_8_n64), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_8_n50), .Q(
        my_filter_q_reg_chain_9__13_), .QN(
        my_filter_delay_line_delay_chain_8_n65) );
  NAND2_X1 my_filter_delay_line_delay_chain_9_U34 ( .A1(
        my_filter_delay_line_n8), .A2(my_filter_q_reg_chain_9__13_), .ZN(
        my_filter_delay_line_delay_chain_9_n92) );
  OAI21_X1 my_filter_delay_line_delay_chain_9_U33 ( .B1(
        my_filter_delay_line_delay_chain_9_n93), .B2(
        my_filter_delay_line_delay_chain_9_n65), .A(
        my_filter_delay_line_delay_chain_9_n92), .ZN(
        my_filter_delay_line_delay_chain_9_n64) );
  NAND2_X1 my_filter_delay_line_delay_chain_9_U32 ( .A1(
        my_filter_q_reg_chain_9__12_), .A2(
        my_filter_delay_line_delay_chain_9_n48), .ZN(
        my_filter_delay_line_delay_chain_9_n91) );
  OAI21_X1 my_filter_delay_line_delay_chain_9_U31 ( .B1(
        my_filter_delay_line_delay_chain_9_n93), .B2(
        my_filter_delay_line_delay_chain_9_n66), .A(
        my_filter_delay_line_delay_chain_9_n91), .ZN(
        my_filter_delay_line_delay_chain_9_n63) );
  NAND2_X1 my_filter_delay_line_delay_chain_9_U30 ( .A1(
        my_filter_q_reg_chain_9__11_), .A2(
        my_filter_delay_line_delay_chain_9_n48), .ZN(
        my_filter_delay_line_delay_chain_9_n90) );
  OAI21_X1 my_filter_delay_line_delay_chain_9_U29 ( .B1(
        my_filter_delay_line_delay_chain_9_n93), .B2(
        my_filter_delay_line_delay_chain_9_n67), .A(
        my_filter_delay_line_delay_chain_9_n90), .ZN(
        my_filter_delay_line_delay_chain_9_n62) );
  NAND2_X1 my_filter_delay_line_delay_chain_9_U28 ( .A1(
        my_filter_q_reg_chain_9__10_), .A2(
        my_filter_delay_line_delay_chain_9_n48), .ZN(
        my_filter_delay_line_delay_chain_9_n89) );
  OAI21_X1 my_filter_delay_line_delay_chain_9_U27 ( .B1(
        my_filter_delay_line_delay_chain_9_n93), .B2(
        my_filter_delay_line_delay_chain_9_n68), .A(
        my_filter_delay_line_delay_chain_9_n89), .ZN(
        my_filter_delay_line_delay_chain_9_n61) );
  NAND2_X1 my_filter_delay_line_delay_chain_9_U26 ( .A1(
        my_filter_q_reg_chain_9__9_), .A2(
        my_filter_delay_line_delay_chain_9_n48), .ZN(
        my_filter_delay_line_delay_chain_9_n88) );
  OAI21_X1 my_filter_delay_line_delay_chain_9_U25 ( .B1(
        my_filter_delay_line_delay_chain_9_n93), .B2(
        my_filter_delay_line_delay_chain_9_n69), .A(
        my_filter_delay_line_delay_chain_9_n88), .ZN(
        my_filter_delay_line_delay_chain_9_n60) );
  NAND2_X1 my_filter_delay_line_delay_chain_9_U24 ( .A1(
        my_filter_q_reg_chain_9__8_), .A2(
        my_filter_delay_line_delay_chain_9_n48), .ZN(
        my_filter_delay_line_delay_chain_9_n87) );
  OAI21_X1 my_filter_delay_line_delay_chain_9_U23 ( .B1(
        my_filter_delay_line_delay_chain_9_n93), .B2(
        my_filter_delay_line_delay_chain_9_n70), .A(
        my_filter_delay_line_delay_chain_9_n87), .ZN(
        my_filter_delay_line_delay_chain_9_n59) );
  NAND2_X1 my_filter_delay_line_delay_chain_9_U22 ( .A1(
        my_filter_q_reg_chain_9__7_), .A2(
        my_filter_delay_line_delay_chain_9_n48), .ZN(
        my_filter_delay_line_delay_chain_9_n86) );
  OAI21_X1 my_filter_delay_line_delay_chain_9_U21 ( .B1(
        my_filter_delay_line_delay_chain_9_n93), .B2(
        my_filter_delay_line_delay_chain_9_n71), .A(
        my_filter_delay_line_delay_chain_9_n86), .ZN(
        my_filter_delay_line_delay_chain_9_n58) );
  NAND2_X1 my_filter_delay_line_delay_chain_9_U20 ( .A1(
        my_filter_q_reg_chain_9__6_), .A2(
        my_filter_delay_line_delay_chain_9_n48), .ZN(
        my_filter_delay_line_delay_chain_9_n85) );
  OAI21_X1 my_filter_delay_line_delay_chain_9_U19 ( .B1(
        my_filter_delay_line_delay_chain_9_n93), .B2(
        my_filter_delay_line_delay_chain_9_n72), .A(
        my_filter_delay_line_delay_chain_9_n85), .ZN(
        my_filter_delay_line_delay_chain_9_n57) );
  NAND2_X1 my_filter_delay_line_delay_chain_9_U18 ( .A1(
        my_filter_q_reg_chain_9__5_), .A2(
        my_filter_delay_line_delay_chain_9_n48), .ZN(
        my_filter_delay_line_delay_chain_9_n84) );
  OAI21_X1 my_filter_delay_line_delay_chain_9_U17 ( .B1(
        my_filter_delay_line_delay_chain_9_n93), .B2(
        my_filter_delay_line_delay_chain_9_n73), .A(
        my_filter_delay_line_delay_chain_9_n84), .ZN(
        my_filter_delay_line_delay_chain_9_n56) );
  NAND2_X1 my_filter_delay_line_delay_chain_9_U16 ( .A1(
        my_filter_q_reg_chain_9__4_), .A2(
        my_filter_delay_line_delay_chain_9_n48), .ZN(
        my_filter_delay_line_delay_chain_9_n83) );
  OAI21_X1 my_filter_delay_line_delay_chain_9_U15 ( .B1(
        my_filter_delay_line_delay_chain_9_n93), .B2(
        my_filter_delay_line_delay_chain_9_n74), .A(
        my_filter_delay_line_delay_chain_9_n83), .ZN(
        my_filter_delay_line_delay_chain_9_n55) );
  NAND2_X1 my_filter_delay_line_delay_chain_9_U14 ( .A1(
        my_filter_q_reg_chain_9__3_), .A2(
        my_filter_delay_line_delay_chain_9_n48), .ZN(
        my_filter_delay_line_delay_chain_9_n82) );
  OAI21_X1 my_filter_delay_line_delay_chain_9_U13 ( .B1(
        my_filter_delay_line_delay_chain_9_n93), .B2(
        my_filter_delay_line_delay_chain_9_n75), .A(
        my_filter_delay_line_delay_chain_9_n82), .ZN(
        my_filter_delay_line_delay_chain_9_n54) );
  NAND2_X1 my_filter_delay_line_delay_chain_9_U12 ( .A1(
        my_filter_q_reg_chain_9__2_), .A2(
        my_filter_delay_line_delay_chain_9_n48), .ZN(
        my_filter_delay_line_delay_chain_9_n81) );
  OAI21_X1 my_filter_delay_line_delay_chain_9_U11 ( .B1(
        my_filter_delay_line_delay_chain_9_n93), .B2(
        my_filter_delay_line_delay_chain_9_n76), .A(
        my_filter_delay_line_delay_chain_9_n81), .ZN(
        my_filter_delay_line_delay_chain_9_n53) );
  NAND2_X1 my_filter_delay_line_delay_chain_9_U10 ( .A1(
        my_filter_q_reg_chain_9__1_), .A2(
        my_filter_delay_line_delay_chain_9_n48), .ZN(
        my_filter_delay_line_delay_chain_9_n80) );
  OAI21_X1 my_filter_delay_line_delay_chain_9_U9 ( .B1(
        my_filter_delay_line_delay_chain_9_n93), .B2(
        my_filter_delay_line_delay_chain_9_n77), .A(
        my_filter_delay_line_delay_chain_9_n80), .ZN(
        my_filter_delay_line_delay_chain_9_n52) );
  NAND2_X1 my_filter_delay_line_delay_chain_9_U8 ( .A1(
        my_filter_q_reg_chain_9__0_), .A2(
        my_filter_delay_line_delay_chain_9_n48), .ZN(
        my_filter_delay_line_delay_chain_9_n79) );
  OAI21_X1 my_filter_delay_line_delay_chain_9_U7 ( .B1(
        my_filter_delay_line_delay_chain_9_n93), .B2(
        my_filter_delay_line_delay_chain_9_n78), .A(
        my_filter_delay_line_delay_chain_9_n79), .ZN(
        my_filter_delay_line_delay_chain_9_n51) );
  INV_X1 my_filter_delay_line_delay_chain_9_U6 ( .A(my_filter_delay_line_n8), 
        .ZN(my_filter_delay_line_delay_chain_9_n49) );
  INV_X1 my_filter_delay_line_delay_chain_9_U5 ( .A(
        my_filter_delay_line_delay_chain_9_n49), .ZN(
        my_filter_delay_line_delay_chain_9_n48) );
  NAND2_X1 my_filter_delay_line_delay_chain_9_U4 ( .A1(
        my_filter_delay_line_delay_chain_9_n50), .A2(
        my_filter_delay_line_delay_chain_9_n49), .ZN(
        my_filter_delay_line_delay_chain_9_n93) );
  BUF_X1 my_filter_delay_line_delay_chain_9_U3 ( .A(my_filter_delay_line_n15), 
        .Z(my_filter_delay_line_delay_chain_9_n50) );
  DFFR_X1 my_filter_delay_line_delay_chain_9_q_reg_0_ ( .D(
        my_filter_delay_line_delay_chain_9_n51), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_9_n50), .Q(
        my_filter_q_reg_chain_10__0_), .QN(
        my_filter_delay_line_delay_chain_9_n78) );
  DFFR_X1 my_filter_delay_line_delay_chain_9_q_reg_1_ ( .D(
        my_filter_delay_line_delay_chain_9_n52), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_9_n50), .Q(
        my_filter_q_reg_chain_10__1_), .QN(
        my_filter_delay_line_delay_chain_9_n77) );
  DFFR_X1 my_filter_delay_line_delay_chain_9_q_reg_2_ ( .D(
        my_filter_delay_line_delay_chain_9_n53), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_9_n50), .Q(
        my_filter_q_reg_chain_10__2_), .QN(
        my_filter_delay_line_delay_chain_9_n76) );
  DFFR_X1 my_filter_delay_line_delay_chain_9_q_reg_3_ ( .D(
        my_filter_delay_line_delay_chain_9_n54), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_9_n50), .Q(
        my_filter_q_reg_chain_10__3_), .QN(
        my_filter_delay_line_delay_chain_9_n75) );
  DFFR_X1 my_filter_delay_line_delay_chain_9_q_reg_4_ ( .D(
        my_filter_delay_line_delay_chain_9_n55), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_9_n50), .Q(
        my_filter_q_reg_chain_10__4_), .QN(
        my_filter_delay_line_delay_chain_9_n74) );
  DFFR_X1 my_filter_delay_line_delay_chain_9_q_reg_5_ ( .D(
        my_filter_delay_line_delay_chain_9_n56), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_9_n50), .Q(
        my_filter_q_reg_chain_10__5_), .QN(
        my_filter_delay_line_delay_chain_9_n73) );
  DFFR_X1 my_filter_delay_line_delay_chain_9_q_reg_6_ ( .D(
        my_filter_delay_line_delay_chain_9_n57), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_9_n50), .Q(
        my_filter_q_reg_chain_10__6_), .QN(
        my_filter_delay_line_delay_chain_9_n72) );
  DFFR_X1 my_filter_delay_line_delay_chain_9_q_reg_7_ ( .D(
        my_filter_delay_line_delay_chain_9_n58), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_9_n50), .Q(
        my_filter_q_reg_chain_10__7_), .QN(
        my_filter_delay_line_delay_chain_9_n71) );
  DFFR_X1 my_filter_delay_line_delay_chain_9_q_reg_8_ ( .D(
        my_filter_delay_line_delay_chain_9_n59), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_9_n50), .Q(
        my_filter_q_reg_chain_10__8_), .QN(
        my_filter_delay_line_delay_chain_9_n70) );
  DFFR_X1 my_filter_delay_line_delay_chain_9_q_reg_9_ ( .D(
        my_filter_delay_line_delay_chain_9_n60), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_9_n50), .Q(
        my_filter_q_reg_chain_10__9_), .QN(
        my_filter_delay_line_delay_chain_9_n69) );
  DFFR_X1 my_filter_delay_line_delay_chain_9_q_reg_10_ ( .D(
        my_filter_delay_line_delay_chain_9_n61), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_9_n50), .Q(
        my_filter_q_reg_chain_10__10_), .QN(
        my_filter_delay_line_delay_chain_9_n68) );
  DFFR_X1 my_filter_delay_line_delay_chain_9_q_reg_11_ ( .D(
        my_filter_delay_line_delay_chain_9_n62), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_9_n50), .Q(
        my_filter_q_reg_chain_10__11_), .QN(
        my_filter_delay_line_delay_chain_9_n67) );
  DFFR_X1 my_filter_delay_line_delay_chain_9_q_reg_12_ ( .D(
        my_filter_delay_line_delay_chain_9_n63), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_9_n50), .Q(
        my_filter_q_reg_chain_10__12_), .QN(
        my_filter_delay_line_delay_chain_9_n66) );
  DFFR_X1 my_filter_delay_line_delay_chain_9_q_reg_13_ ( .D(
        my_filter_delay_line_delay_chain_9_n64), .CK(clk), .RN(
        my_filter_delay_line_delay_chain_9_n50), .Q(
        my_filter_q_reg_chain_10__13_), .QN(
        my_filter_delay_line_delay_chain_9_n65) );
  NOR2_X1 my_filter_first_coeff_mult_21_U276 ( .A1(
        my_filter_first_coeff_mult_21_n87), .A2(
        my_filter_first_coeff_mult_21_n101), .ZN(
        my_filter_first_coeff_mult_21_ab_12__12_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U275 ( .A1(my_filter_q_reg_samp_11_), 
        .A2(my_filter_first_coeff_mult_21_n86), .ZN(
        my_filter_first_coeff_mult_21_ab_11__13_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U274 ( .A1(
        my_filter_first_coeff_mult_21_n87), .A2(
        my_filter_first_coeff_mult_21_n102), .ZN(
        my_filter_first_coeff_mult_21_ab_11__12_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U273 ( .A1(my_filter_q_reg_samp_10_), 
        .A2(my_filter_first_coeff_mult_21_n86), .ZN(
        my_filter_first_coeff_mult_21_ab_10__13_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U272 ( .A1(
        my_filter_first_coeff_mult_21_n87), .A2(
        my_filter_first_coeff_mult_21_n103), .ZN(
        my_filter_first_coeff_mult_21_ab_10__12_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U271 ( .A1(my_filter_q_reg_samp_9_), 
        .A2(my_filter_first_coeff_mult_21_n86), .ZN(
        my_filter_first_coeff_mult_21_ab_9__13_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U270 ( .A1(my_filter_q_reg_samp_8_), 
        .A2(my_filter_first_coeff_mult_21_n86), .ZN(
        my_filter_first_coeff_mult_21_ab_8__13_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U269 ( .A1(
        my_filter_first_coeff_mult_21_n104), .A2(
        my_filter_first_coeff_mult_21_n87), .ZN(
        my_filter_first_coeff_mult_21_ab_9__12_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U268 ( .A1(my_filter_q_reg_coeff[150]), 
        .A2(my_filter_first_coeff_mult_21_n100), .ZN(
        my_filter_first_coeff_mult_21_ab_13__10_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U267 ( .A1(my_filter_q_reg_coeff[151]), 
        .A2(my_filter_first_coeff_mult_21_n100), .ZN(
        my_filter_first_coeff_mult_21_ab_13__11_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U266 ( .A1(my_filter_q_reg_coeff[149]), 
        .A2(my_filter_first_coeff_mult_21_n100), .ZN(
        my_filter_first_coeff_mult_21_ab_13__9_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U265 ( .A1(my_filter_q_reg_coeff[152]), 
        .A2(my_filter_first_coeff_mult_21_n100), .ZN(
        my_filter_first_coeff_mult_21_ab_13__12_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U264 ( .A1(my_filter_q_reg_samp_12_), 
        .A2(my_filter_first_coeff_mult_21_n86), .ZN(
        my_filter_first_coeff_mult_21_ab_12__13_) );
  INV_X1 my_filter_first_coeff_mult_21_U263 ( .A(my_filter_q_reg_samp_9_), 
        .ZN(my_filter_first_coeff_mult_21_n104) );
  INV_X1 my_filter_first_coeff_mult_21_U262 ( .A(my_filter_q_reg_samp_12_), 
        .ZN(my_filter_first_coeff_mult_21_n101) );
  INV_X1 my_filter_first_coeff_mult_21_U261 ( .A(my_filter_q_reg_samp_11_), 
        .ZN(my_filter_first_coeff_mult_21_n102) );
  INV_X1 my_filter_first_coeff_mult_21_U260 ( .A(my_filter_q_reg_samp_10_), 
        .ZN(my_filter_first_coeff_mult_21_n103) );
  INV_X1 my_filter_first_coeff_mult_21_U259 ( .A(my_filter_q_reg_samp_8_), 
        .ZN(my_filter_first_coeff_mult_21_n105) );
  INV_X1 my_filter_first_coeff_mult_21_U258 ( .A(my_filter_q_reg_samp_13_), 
        .ZN(my_filter_first_coeff_mult_21_n100) );
  AND2_X1 my_filter_first_coeff_mult_21_U257 ( .A1(
        my_filter_first_coeff_mult_21_ab_0__13_), .A2(
        my_filter_first_coeff_mult_21_ab_1__12_), .ZN(
        my_filter_first_coeff_mult_21_n15) );
  NOR2_X1 my_filter_first_coeff_mult_21_U256 ( .A1(
        my_filter_first_coeff_mult_21_n87), .A2(
        my_filter_first_coeff_mult_21_n111), .ZN(
        my_filter_first_coeff_mult_21_ab_2__12_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U255 ( .A1(my_filter_q_reg_samp_1_), 
        .A2(my_filter_first_coeff_mult_21_n86), .ZN(
        my_filter_first_coeff_mult_21_ab_1__13_) );
  AND3_X1 my_filter_first_coeff_mult_21_U254 ( .A1(
        my_filter_first_coeff_mult_21_ab_1__1_), .A2(
        my_filter_q_reg_coeff[140]), .A3(my_filter_q_reg_samp_0_), .ZN(
        my_filter_first_coeff_mult_21_CARRYB_1__0_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U253 ( .A1(
        my_filter_first_coeff_mult_21_n99), .A2(
        my_filter_first_coeff_mult_21_n101), .ZN(
        my_filter_first_coeff_mult_21_ab_12__0_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U252 ( .A1(my_filter_q_reg_coeff[140]), 
        .A2(my_filter_first_coeff_mult_21_n100), .ZN(
        my_filter_first_coeff_mult_21_ab_13__0_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U251 ( .A1(
        my_filter_first_coeff_mult_21_n87), .A2(
        my_filter_first_coeff_mult_21_n105), .ZN(
        my_filter_first_coeff_mult_21_ab_8__12_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U250 ( .A1(my_filter_q_reg_samp_7_), 
        .A2(my_filter_first_coeff_mult_21_n86), .ZN(
        my_filter_first_coeff_mult_21_ab_7__13_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U249 ( .A1(
        my_filter_first_coeff_mult_21_n87), .A2(
        my_filter_first_coeff_mult_21_n106), .ZN(
        my_filter_first_coeff_mult_21_ab_7__12_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U248 ( .A1(my_filter_q_reg_samp_6_), 
        .A2(my_filter_first_coeff_mult_21_n86), .ZN(
        my_filter_first_coeff_mult_21_ab_6__13_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U247 ( .A1(
        my_filter_first_coeff_mult_21_n87), .A2(
        my_filter_first_coeff_mult_21_n107), .ZN(
        my_filter_first_coeff_mult_21_ab_6__12_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U246 ( .A1(my_filter_q_reg_samp_5_), 
        .A2(my_filter_first_coeff_mult_21_n86), .ZN(
        my_filter_first_coeff_mult_21_ab_5__13_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U245 ( .A1(
        my_filter_first_coeff_mult_21_n87), .A2(
        my_filter_first_coeff_mult_21_n108), .ZN(
        my_filter_first_coeff_mult_21_ab_5__12_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U244 ( .A1(my_filter_q_reg_samp_4_), 
        .A2(my_filter_first_coeff_mult_21_n86), .ZN(
        my_filter_first_coeff_mult_21_ab_4__13_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U243 ( .A1(
        my_filter_first_coeff_mult_21_n87), .A2(
        my_filter_first_coeff_mult_21_n109), .ZN(
        my_filter_first_coeff_mult_21_ab_4__12_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U242 ( .A1(my_filter_q_reg_samp_3_), 
        .A2(my_filter_first_coeff_mult_21_n86), .ZN(
        my_filter_first_coeff_mult_21_ab_3__13_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U241 ( .A1(
        my_filter_first_coeff_mult_21_n87), .A2(
        my_filter_first_coeff_mult_21_n110), .ZN(
        my_filter_first_coeff_mult_21_ab_3__12_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U240 ( .A1(my_filter_q_reg_samp_2_), 
        .A2(my_filter_first_coeff_mult_21_n86), .ZN(
        my_filter_first_coeff_mult_21_ab_2__13_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U239 ( .A1(my_filter_q_reg_coeff[148]), 
        .A2(my_filter_first_coeff_mult_21_n100), .ZN(
        my_filter_first_coeff_mult_21_ab_13__8_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U238 ( .A1(my_filter_q_reg_coeff[146]), 
        .A2(my_filter_first_coeff_mult_21_n100), .ZN(
        my_filter_first_coeff_mult_21_ab_13__6_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U237 ( .A1(my_filter_q_reg_coeff[147]), 
        .A2(my_filter_first_coeff_mult_21_n100), .ZN(
        my_filter_first_coeff_mult_21_ab_13__7_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U236 ( .A1(my_filter_q_reg_coeff[144]), 
        .A2(my_filter_first_coeff_mult_21_n100), .ZN(
        my_filter_first_coeff_mult_21_ab_13__4_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U235 ( .A1(my_filter_q_reg_coeff[145]), 
        .A2(my_filter_first_coeff_mult_21_n100), .ZN(
        my_filter_first_coeff_mult_21_ab_13__5_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U234 ( .A1(my_filter_q_reg_coeff[142]), 
        .A2(my_filter_first_coeff_mult_21_n100), .ZN(
        my_filter_first_coeff_mult_21_ab_13__2_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U233 ( .A1(my_filter_q_reg_coeff[143]), 
        .A2(my_filter_first_coeff_mult_21_n100), .ZN(
        my_filter_first_coeff_mult_21_ab_13__3_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U232 ( .A1(my_filter_q_reg_coeff[141]), 
        .A2(my_filter_first_coeff_mult_21_n100), .ZN(
        my_filter_first_coeff_mult_21_ab_13__1_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U231 ( .A1(my_filter_q_reg_samp_0_), 
        .A2(my_filter_first_coeff_mult_21_n86), .ZN(
        my_filter_first_coeff_mult_21_ab_0__13_) );
  INV_X1 my_filter_first_coeff_mult_21_U230 ( .A(my_filter_q_reg_coeff[153]), 
        .ZN(my_filter_first_coeff_mult_21_n86) );
  INV_X1 my_filter_first_coeff_mult_21_U229 ( .A(my_filter_q_reg_coeff[140]), 
        .ZN(my_filter_first_coeff_mult_21_n99) );
  INV_X1 my_filter_first_coeff_mult_21_U228 ( .A(my_filter_q_reg_samp_0_), 
        .ZN(my_filter_first_coeff_mult_21_n113) );
  INV_X1 my_filter_first_coeff_mult_21_U227 ( .A(my_filter_q_reg_coeff[141]), 
        .ZN(my_filter_first_coeff_mult_21_n98) );
  INV_X1 my_filter_first_coeff_mult_21_U226 ( .A(my_filter_q_reg_samp_1_), 
        .ZN(my_filter_first_coeff_mult_21_n112) );
  INV_X1 my_filter_first_coeff_mult_21_U225 ( .A(my_filter_q_reg_coeff[152]), 
        .ZN(my_filter_first_coeff_mult_21_n87) );
  INV_X1 my_filter_first_coeff_mult_21_U224 ( .A(my_filter_q_reg_coeff[150]), 
        .ZN(my_filter_first_coeff_mult_21_n89) );
  INV_X1 my_filter_first_coeff_mult_21_U223 ( .A(my_filter_q_reg_coeff[151]), 
        .ZN(my_filter_first_coeff_mult_21_n88) );
  INV_X1 my_filter_first_coeff_mult_21_U222 ( .A(my_filter_q_reg_coeff[148]), 
        .ZN(my_filter_first_coeff_mult_21_n91) );
  INV_X1 my_filter_first_coeff_mult_21_U221 ( .A(my_filter_q_reg_coeff[149]), 
        .ZN(my_filter_first_coeff_mult_21_n90) );
  INV_X1 my_filter_first_coeff_mult_21_U220 ( .A(my_filter_q_reg_coeff[146]), 
        .ZN(my_filter_first_coeff_mult_21_n93) );
  INV_X1 my_filter_first_coeff_mult_21_U219 ( .A(my_filter_q_reg_coeff[147]), 
        .ZN(my_filter_first_coeff_mult_21_n92) );
  INV_X1 my_filter_first_coeff_mult_21_U218 ( .A(my_filter_q_reg_coeff[142]), 
        .ZN(my_filter_first_coeff_mult_21_n97) );
  INV_X1 my_filter_first_coeff_mult_21_U217 ( .A(my_filter_q_reg_coeff[143]), 
        .ZN(my_filter_first_coeff_mult_21_n96) );
  INV_X1 my_filter_first_coeff_mult_21_U216 ( .A(my_filter_q_reg_coeff[144]), 
        .ZN(my_filter_first_coeff_mult_21_n95) );
  INV_X1 my_filter_first_coeff_mult_21_U215 ( .A(my_filter_q_reg_coeff[145]), 
        .ZN(my_filter_first_coeff_mult_21_n94) );
  INV_X1 my_filter_first_coeff_mult_21_U214 ( .A(my_filter_q_reg_samp_7_), 
        .ZN(my_filter_first_coeff_mult_21_n106) );
  INV_X1 my_filter_first_coeff_mult_21_U213 ( .A(my_filter_q_reg_samp_6_), 
        .ZN(my_filter_first_coeff_mult_21_n107) );
  INV_X1 my_filter_first_coeff_mult_21_U212 ( .A(my_filter_q_reg_samp_5_), 
        .ZN(my_filter_first_coeff_mult_21_n108) );
  INV_X1 my_filter_first_coeff_mult_21_U211 ( .A(my_filter_q_reg_samp_4_), 
        .ZN(my_filter_first_coeff_mult_21_n109) );
  INV_X1 my_filter_first_coeff_mult_21_U210 ( .A(my_filter_q_reg_samp_2_), 
        .ZN(my_filter_first_coeff_mult_21_n111) );
  INV_X1 my_filter_first_coeff_mult_21_U209 ( .A(my_filter_q_reg_samp_3_), 
        .ZN(my_filter_first_coeff_mult_21_n110) );
  AND2_X1 my_filter_first_coeff_mult_21_U208 ( .A1(
        my_filter_first_coeff_mult_21_CARRYB_13__12_), .A2(
        my_filter_first_coeff_mult_21_SUMB_13__13_), .ZN(
        my_filter_first_coeff_mult_21_n3) );
  NOR2_X1 my_filter_first_coeff_mult_21_U207 ( .A1(
        my_filter_first_coeff_mult_21_n86), .A2(
        my_filter_first_coeff_mult_21_n100), .ZN(
        my_filter_first_coeff_mult_21_ab_13__13_) );
  AND2_X1 my_filter_first_coeff_mult_21_U206 ( .A1(
        my_filter_first_coeff_mult_21_CARRYB_13__11_), .A2(
        my_filter_first_coeff_mult_21_SUMB_13__12_), .ZN(
        my_filter_first_coeff_mult_21_n27) );
  AND2_X1 my_filter_first_coeff_mult_21_U205 ( .A1(
        my_filter_first_coeff_mult_21_CARRYB_13__9_), .A2(
        my_filter_first_coeff_mult_21_SUMB_13__10_), .ZN(
        my_filter_first_coeff_mult_21_n52) );
  AND2_X1 my_filter_first_coeff_mult_21_U204 ( .A1(
        my_filter_first_coeff_mult_21_CARRYB_13__7_), .A2(
        my_filter_first_coeff_mult_21_SUMB_13__8_), .ZN(
        my_filter_first_coeff_mult_21_n51) );
  AND2_X1 my_filter_first_coeff_mult_21_U203 ( .A1(
        my_filter_first_coeff_mult_21_CARRYB_13__10_), .A2(
        my_filter_first_coeff_mult_21_SUMB_13__11_), .ZN(
        my_filter_first_coeff_mult_21_n48) );
  AND2_X1 my_filter_first_coeff_mult_21_U202 ( .A1(
        my_filter_first_coeff_mult_21_CARRYB_13__8_), .A2(
        my_filter_first_coeff_mult_21_SUMB_13__9_), .ZN(
        my_filter_first_coeff_mult_21_n49) );
  AND2_X1 my_filter_first_coeff_mult_21_U201 ( .A1(
        my_filter_first_coeff_mult_21_CARRYB_13__6_), .A2(
        my_filter_first_coeff_mult_21_SUMB_13__7_), .ZN(
        my_filter_first_coeff_mult_21_n41) );
  NOR2_X1 my_filter_first_coeff_mult_21_U200 ( .A1(
        my_filter_first_coeff_mult_21_n88), .A2(
        my_filter_first_coeff_mult_21_n101), .ZN(
        my_filter_first_coeff_mult_21_ab_12__11_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U199 ( .A1(
        my_filter_first_coeff_mult_21_n89), .A2(
        my_filter_first_coeff_mult_21_n101), .ZN(
        my_filter_first_coeff_mult_21_ab_12__10_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U198 ( .A1(
        my_filter_first_coeff_mult_21_n88), .A2(
        my_filter_first_coeff_mult_21_n102), .ZN(
        my_filter_first_coeff_mult_21_ab_11__11_) );
  AND2_X1 my_filter_first_coeff_mult_21_U197 ( .A1(
        my_filter_first_coeff_mult_21_CARRYB_13__5_), .A2(
        my_filter_first_coeff_mult_21_SUMB_13__6_), .ZN(
        my_filter_first_coeff_mult_21_n43) );
  AND2_X1 my_filter_first_coeff_mult_21_U196 ( .A1(
        my_filter_first_coeff_mult_21_CARRYB_13__3_), .A2(
        my_filter_first_coeff_mult_21_SUMB_13__4_), .ZN(
        my_filter_first_coeff_mult_21_n34) );
  AND2_X1 my_filter_first_coeff_mult_21_U195 ( .A1(
        my_filter_first_coeff_mult_21_CARRYB_13__1_), .A2(
        my_filter_first_coeff_mult_21_SUMB_13__2_), .ZN(
        my_filter_first_coeff_mult_21_n42) );
  AND2_X1 my_filter_first_coeff_mult_21_U194 ( .A1(
        my_filter_first_coeff_mult_21_CARRYB_13__4_), .A2(
        my_filter_first_coeff_mult_21_SUMB_13__5_), .ZN(
        my_filter_first_coeff_mult_21_n40) );
  AND2_X1 my_filter_first_coeff_mult_21_U193 ( .A1(
        my_filter_first_coeff_mult_21_CARRYB_13__2_), .A2(
        my_filter_first_coeff_mult_21_SUMB_13__3_), .ZN(
        my_filter_first_coeff_mult_21_n39) );
  AND2_X1 my_filter_first_coeff_mult_21_U192 ( .A1(
        my_filter_first_coeff_mult_21_CARRYB_13__0_), .A2(
        my_filter_first_coeff_mult_21_SUMB_13__1_), .ZN(
        my_filter_first_coeff_mult_21_n38) );
  NOR2_X1 my_filter_first_coeff_mult_21_U191 ( .A1(
        my_filter_first_coeff_mult_21_n99), .A2(
        my_filter_first_coeff_mult_21_n103), .ZN(
        my_filter_first_coeff_mult_21_ab_10__0_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U190 ( .A1(
        my_filter_first_coeff_mult_21_n99), .A2(
        my_filter_first_coeff_mult_21_n102), .ZN(
        my_filter_first_coeff_mult_21_ab_11__0_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U189 ( .A1(
        my_filter_first_coeff_mult_21_n98), .A2(
        my_filter_first_coeff_mult_21_n102), .ZN(
        my_filter_first_coeff_mult_21_ab_11__1_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U188 ( .A1(
        my_filter_first_coeff_mult_21_n98), .A2(
        my_filter_first_coeff_mult_21_n103), .ZN(
        my_filter_first_coeff_mult_21_ab_10__1_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U187 ( .A1(
        my_filter_first_coeff_mult_21_n99), .A2(
        my_filter_first_coeff_mult_21_n105), .ZN(
        my_filter_first_coeff_mult_21_ab_8__0_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U186 ( .A1(
        my_filter_first_coeff_mult_21_n104), .A2(
        my_filter_first_coeff_mult_21_n99), .ZN(
        my_filter_first_coeff_mult_21_ab_9__0_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U185 ( .A1(
        my_filter_first_coeff_mult_21_n104), .A2(
        my_filter_first_coeff_mult_21_n98), .ZN(
        my_filter_first_coeff_mult_21_ab_9__1_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U184 ( .A1(
        my_filter_first_coeff_mult_21_n104), .A2(
        my_filter_first_coeff_mult_21_n97), .ZN(
        my_filter_first_coeff_mult_21_ab_9__2_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U183 ( .A1(
        my_filter_first_coeff_mult_21_n104), .A2(
        my_filter_first_coeff_mult_21_n96), .ZN(
        my_filter_first_coeff_mult_21_ab_9__3_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U182 ( .A1(
        my_filter_first_coeff_mult_21_n98), .A2(
        my_filter_first_coeff_mult_21_n105), .ZN(
        my_filter_first_coeff_mult_21_ab_8__1_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U181 ( .A1(
        my_filter_first_coeff_mult_21_n96), .A2(
        my_filter_first_coeff_mult_21_n105), .ZN(
        my_filter_first_coeff_mult_21_ab_8__3_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U180 ( .A1(
        my_filter_first_coeff_mult_21_n99), .A2(
        my_filter_first_coeff_mult_21_n107), .ZN(
        my_filter_first_coeff_mult_21_ab_6__0_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U179 ( .A1(
        my_filter_first_coeff_mult_21_n99), .A2(
        my_filter_first_coeff_mult_21_n106), .ZN(
        my_filter_first_coeff_mult_21_ab_7__0_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U178 ( .A1(
        my_filter_first_coeff_mult_21_n98), .A2(
        my_filter_first_coeff_mult_21_n106), .ZN(
        my_filter_first_coeff_mult_21_ab_7__1_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U177 ( .A1(
        my_filter_first_coeff_mult_21_n97), .A2(
        my_filter_first_coeff_mult_21_n106), .ZN(
        my_filter_first_coeff_mult_21_ab_7__2_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U176 ( .A1(
        my_filter_first_coeff_mult_21_n96), .A2(
        my_filter_first_coeff_mult_21_n106), .ZN(
        my_filter_first_coeff_mult_21_ab_7__3_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U175 ( .A1(
        my_filter_first_coeff_mult_21_n95), .A2(
        my_filter_first_coeff_mult_21_n106), .ZN(
        my_filter_first_coeff_mult_21_ab_7__4_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U174 ( .A1(
        my_filter_first_coeff_mult_21_n94), .A2(
        my_filter_first_coeff_mult_21_n106), .ZN(
        my_filter_first_coeff_mult_21_ab_7__5_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U173 ( .A1(
        my_filter_first_coeff_mult_21_n98), .A2(
        my_filter_first_coeff_mult_21_n107), .ZN(
        my_filter_first_coeff_mult_21_ab_6__1_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U172 ( .A1(
        my_filter_first_coeff_mult_21_n96), .A2(
        my_filter_first_coeff_mult_21_n107), .ZN(
        my_filter_first_coeff_mult_21_ab_6__3_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U171 ( .A1(
        my_filter_first_coeff_mult_21_n94), .A2(
        my_filter_first_coeff_mult_21_n107), .ZN(
        my_filter_first_coeff_mult_21_ab_6__5_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U170 ( .A1(
        my_filter_first_coeff_mult_21_n99), .A2(
        my_filter_first_coeff_mult_21_n109), .ZN(
        my_filter_first_coeff_mult_21_ab_4__0_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U169 ( .A1(
        my_filter_first_coeff_mult_21_n99), .A2(
        my_filter_first_coeff_mult_21_n108), .ZN(
        my_filter_first_coeff_mult_21_ab_5__0_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U168 ( .A1(
        my_filter_first_coeff_mult_21_n98), .A2(
        my_filter_first_coeff_mult_21_n108), .ZN(
        my_filter_first_coeff_mult_21_ab_5__1_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U167 ( .A1(
        my_filter_first_coeff_mult_21_n97), .A2(
        my_filter_first_coeff_mult_21_n108), .ZN(
        my_filter_first_coeff_mult_21_ab_5__2_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U166 ( .A1(
        my_filter_first_coeff_mult_21_n96), .A2(
        my_filter_first_coeff_mult_21_n108), .ZN(
        my_filter_first_coeff_mult_21_ab_5__3_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U165 ( .A1(
        my_filter_first_coeff_mult_21_n95), .A2(
        my_filter_first_coeff_mult_21_n108), .ZN(
        my_filter_first_coeff_mult_21_ab_5__4_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U164 ( .A1(
        my_filter_first_coeff_mult_21_n94), .A2(
        my_filter_first_coeff_mult_21_n108), .ZN(
        my_filter_first_coeff_mult_21_ab_5__5_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U163 ( .A1(
        my_filter_first_coeff_mult_21_n93), .A2(
        my_filter_first_coeff_mult_21_n108), .ZN(
        my_filter_first_coeff_mult_21_ab_5__6_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U162 ( .A1(
        my_filter_first_coeff_mult_21_n92), .A2(
        my_filter_first_coeff_mult_21_n108), .ZN(
        my_filter_first_coeff_mult_21_ab_5__7_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U161 ( .A1(
        my_filter_first_coeff_mult_21_n98), .A2(
        my_filter_first_coeff_mult_21_n109), .ZN(
        my_filter_first_coeff_mult_21_ab_4__1_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U160 ( .A1(
        my_filter_first_coeff_mult_21_n96), .A2(
        my_filter_first_coeff_mult_21_n109), .ZN(
        my_filter_first_coeff_mult_21_ab_4__3_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U159 ( .A1(
        my_filter_first_coeff_mult_21_n94), .A2(
        my_filter_first_coeff_mult_21_n109), .ZN(
        my_filter_first_coeff_mult_21_ab_4__5_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U158 ( .A1(
        my_filter_first_coeff_mult_21_n99), .A2(
        my_filter_first_coeff_mult_21_n111), .ZN(
        my_filter_first_coeff_mult_21_ab_2__0_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U157 ( .A1(
        my_filter_first_coeff_mult_21_n99), .A2(
        my_filter_first_coeff_mult_21_n110), .ZN(
        my_filter_first_coeff_mult_21_ab_3__0_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U156 ( .A1(
        my_filter_first_coeff_mult_21_n98), .A2(
        my_filter_first_coeff_mult_21_n110), .ZN(
        my_filter_first_coeff_mult_21_ab_3__1_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U155 ( .A1(
        my_filter_first_coeff_mult_21_n97), .A2(
        my_filter_first_coeff_mult_21_n110), .ZN(
        my_filter_first_coeff_mult_21_ab_3__2_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U154 ( .A1(
        my_filter_first_coeff_mult_21_n96), .A2(
        my_filter_first_coeff_mult_21_n110), .ZN(
        my_filter_first_coeff_mult_21_ab_3__3_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U153 ( .A1(
        my_filter_first_coeff_mult_21_n95), .A2(
        my_filter_first_coeff_mult_21_n110), .ZN(
        my_filter_first_coeff_mult_21_ab_3__4_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U152 ( .A1(
        my_filter_first_coeff_mult_21_n94), .A2(
        my_filter_first_coeff_mult_21_n110), .ZN(
        my_filter_first_coeff_mult_21_ab_3__5_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U151 ( .A1(
        my_filter_first_coeff_mult_21_n93), .A2(
        my_filter_first_coeff_mult_21_n110), .ZN(
        my_filter_first_coeff_mult_21_ab_3__6_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U150 ( .A1(
        my_filter_first_coeff_mult_21_n91), .A2(
        my_filter_first_coeff_mult_21_n110), .ZN(
        my_filter_first_coeff_mult_21_ab_3__8_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U149 ( .A1(
        my_filter_first_coeff_mult_21_n90), .A2(
        my_filter_first_coeff_mult_21_n110), .ZN(
        my_filter_first_coeff_mult_21_ab_3__9_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U148 ( .A1(
        my_filter_first_coeff_mult_21_n90), .A2(
        my_filter_first_coeff_mult_21_n101), .ZN(
        my_filter_first_coeff_mult_21_ab_12__9_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U147 ( .A1(
        my_filter_first_coeff_mult_21_n89), .A2(
        my_filter_first_coeff_mult_21_n102), .ZN(
        my_filter_first_coeff_mult_21_ab_11__10_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U146 ( .A1(
        my_filter_first_coeff_mult_21_n92), .A2(
        my_filter_first_coeff_mult_21_n101), .ZN(
        my_filter_first_coeff_mult_21_ab_12__7_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U145 ( .A1(
        my_filter_first_coeff_mult_21_n91), .A2(
        my_filter_first_coeff_mult_21_n101), .ZN(
        my_filter_first_coeff_mult_21_ab_12__8_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U144 ( .A1(
        my_filter_first_coeff_mult_21_n88), .A2(
        my_filter_first_coeff_mult_21_n103), .ZN(
        my_filter_first_coeff_mult_21_ab_10__11_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U143 ( .A1(
        my_filter_first_coeff_mult_21_n91), .A2(
        my_filter_first_coeff_mult_21_n102), .ZN(
        my_filter_first_coeff_mult_21_ab_11__8_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U142 ( .A1(
        my_filter_first_coeff_mult_21_n90), .A2(
        my_filter_first_coeff_mult_21_n102), .ZN(
        my_filter_first_coeff_mult_21_ab_11__9_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U141 ( .A1(
        my_filter_first_coeff_mult_21_n94), .A2(
        my_filter_first_coeff_mult_21_n101), .ZN(
        my_filter_first_coeff_mult_21_ab_12__5_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U140 ( .A1(
        my_filter_first_coeff_mult_21_n93), .A2(
        my_filter_first_coeff_mult_21_n101), .ZN(
        my_filter_first_coeff_mult_21_ab_12__6_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U139 ( .A1(
        my_filter_first_coeff_mult_21_n90), .A2(
        my_filter_first_coeff_mult_21_n103), .ZN(
        my_filter_first_coeff_mult_21_ab_10__9_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U138 ( .A1(
        my_filter_first_coeff_mult_21_n89), .A2(
        my_filter_first_coeff_mult_21_n103), .ZN(
        my_filter_first_coeff_mult_21_ab_10__10_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U137 ( .A1(
        my_filter_first_coeff_mult_21_n93), .A2(
        my_filter_first_coeff_mult_21_n102), .ZN(
        my_filter_first_coeff_mult_21_ab_11__6_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U136 ( .A1(
        my_filter_first_coeff_mult_21_n92), .A2(
        my_filter_first_coeff_mult_21_n102), .ZN(
        my_filter_first_coeff_mult_21_ab_11__7_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U135 ( .A1(
        my_filter_first_coeff_mult_21_n104), .A2(
        my_filter_first_coeff_mult_21_n89), .ZN(
        my_filter_first_coeff_mult_21_ab_9__10_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U134 ( .A1(
        my_filter_first_coeff_mult_21_n104), .A2(
        my_filter_first_coeff_mult_21_n88), .ZN(
        my_filter_first_coeff_mult_21_ab_9__11_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U133 ( .A1(
        my_filter_first_coeff_mult_21_n96), .A2(
        my_filter_first_coeff_mult_21_n101), .ZN(
        my_filter_first_coeff_mult_21_ab_12__3_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U132 ( .A1(
        my_filter_first_coeff_mult_21_n95), .A2(
        my_filter_first_coeff_mult_21_n101), .ZN(
        my_filter_first_coeff_mult_21_ab_12__4_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U131 ( .A1(
        my_filter_first_coeff_mult_21_n92), .A2(
        my_filter_first_coeff_mult_21_n103), .ZN(
        my_filter_first_coeff_mult_21_ab_10__7_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U130 ( .A1(
        my_filter_first_coeff_mult_21_n91), .A2(
        my_filter_first_coeff_mult_21_n103), .ZN(
        my_filter_first_coeff_mult_21_ab_10__8_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U129 ( .A1(
        my_filter_first_coeff_mult_21_n88), .A2(
        my_filter_first_coeff_mult_21_n105), .ZN(
        my_filter_first_coeff_mult_21_ab_8__11_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U128 ( .A1(
        my_filter_first_coeff_mult_21_n97), .A2(
        my_filter_first_coeff_mult_21_n101), .ZN(
        my_filter_first_coeff_mult_21_ab_12__2_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U127 ( .A1(
        my_filter_first_coeff_mult_21_n95), .A2(
        my_filter_first_coeff_mult_21_n102), .ZN(
        my_filter_first_coeff_mult_21_ab_11__4_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U126 ( .A1(
        my_filter_first_coeff_mult_21_n94), .A2(
        my_filter_first_coeff_mult_21_n102), .ZN(
        my_filter_first_coeff_mult_21_ab_11__5_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U125 ( .A1(
        my_filter_first_coeff_mult_21_n104), .A2(
        my_filter_first_coeff_mult_21_n91), .ZN(
        my_filter_first_coeff_mult_21_ab_9__8_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U124 ( .A1(
        my_filter_first_coeff_mult_21_n104), .A2(
        my_filter_first_coeff_mult_21_n90), .ZN(
        my_filter_first_coeff_mult_21_ab_9__9_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U123 ( .A1(
        my_filter_first_coeff_mult_21_n96), .A2(
        my_filter_first_coeff_mult_21_n102), .ZN(
        my_filter_first_coeff_mult_21_ab_11__3_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U122 ( .A1(
        my_filter_first_coeff_mult_21_n98), .A2(
        my_filter_first_coeff_mult_21_n101), .ZN(
        my_filter_first_coeff_mult_21_ab_12__1_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U121 ( .A1(
        my_filter_first_coeff_mult_21_n94), .A2(
        my_filter_first_coeff_mult_21_n103), .ZN(
        my_filter_first_coeff_mult_21_ab_10__5_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U120 ( .A1(
        my_filter_first_coeff_mult_21_n93), .A2(
        my_filter_first_coeff_mult_21_n103), .ZN(
        my_filter_first_coeff_mult_21_ab_10__6_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U119 ( .A1(
        my_filter_first_coeff_mult_21_n90), .A2(
        my_filter_first_coeff_mult_21_n105), .ZN(
        my_filter_first_coeff_mult_21_ab_8__9_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U118 ( .A1(
        my_filter_first_coeff_mult_21_n89), .A2(
        my_filter_first_coeff_mult_21_n105), .ZN(
        my_filter_first_coeff_mult_21_ab_8__10_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U117 ( .A1(
        my_filter_first_coeff_mult_21_n95), .A2(
        my_filter_first_coeff_mult_21_n103), .ZN(
        my_filter_first_coeff_mult_21_ab_10__4_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U116 ( .A1(
        my_filter_first_coeff_mult_21_n97), .A2(
        my_filter_first_coeff_mult_21_n102), .ZN(
        my_filter_first_coeff_mult_21_ab_11__2_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U115 ( .A1(
        my_filter_first_coeff_mult_21_n104), .A2(
        my_filter_first_coeff_mult_21_n93), .ZN(
        my_filter_first_coeff_mult_21_ab_9__6_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U114 ( .A1(
        my_filter_first_coeff_mult_21_n104), .A2(
        my_filter_first_coeff_mult_21_n92), .ZN(
        my_filter_first_coeff_mult_21_ab_9__7_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U113 ( .A1(
        my_filter_first_coeff_mult_21_n89), .A2(
        my_filter_first_coeff_mult_21_n106), .ZN(
        my_filter_first_coeff_mult_21_ab_7__10_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U112 ( .A1(
        my_filter_first_coeff_mult_21_n88), .A2(
        my_filter_first_coeff_mult_21_n106), .ZN(
        my_filter_first_coeff_mult_21_ab_7__11_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U111 ( .A1(
        my_filter_first_coeff_mult_21_n104), .A2(
        my_filter_first_coeff_mult_21_n94), .ZN(
        my_filter_first_coeff_mult_21_ab_9__5_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U110 ( .A1(
        my_filter_first_coeff_mult_21_n97), .A2(
        my_filter_first_coeff_mult_21_n103), .ZN(
        my_filter_first_coeff_mult_21_ab_10__2_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U109 ( .A1(
        my_filter_first_coeff_mult_21_n96), .A2(
        my_filter_first_coeff_mult_21_n103), .ZN(
        my_filter_first_coeff_mult_21_ab_10__3_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U108 ( .A1(
        my_filter_first_coeff_mult_21_n92), .A2(
        my_filter_first_coeff_mult_21_n105), .ZN(
        my_filter_first_coeff_mult_21_ab_8__7_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U107 ( .A1(
        my_filter_first_coeff_mult_21_n91), .A2(
        my_filter_first_coeff_mult_21_n105), .ZN(
        my_filter_first_coeff_mult_21_ab_8__8_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U106 ( .A1(
        my_filter_first_coeff_mult_21_n88), .A2(
        my_filter_first_coeff_mult_21_n107), .ZN(
        my_filter_first_coeff_mult_21_ab_6__11_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U105 ( .A1(
        my_filter_first_coeff_mult_21_n93), .A2(
        my_filter_first_coeff_mult_21_n105), .ZN(
        my_filter_first_coeff_mult_21_ab_8__6_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U104 ( .A1(
        my_filter_first_coeff_mult_21_n104), .A2(
        my_filter_first_coeff_mult_21_n95), .ZN(
        my_filter_first_coeff_mult_21_ab_9__4_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U103 ( .A1(
        my_filter_first_coeff_mult_21_n91), .A2(
        my_filter_first_coeff_mult_21_n106), .ZN(
        my_filter_first_coeff_mult_21_ab_7__8_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U102 ( .A1(
        my_filter_first_coeff_mult_21_n90), .A2(
        my_filter_first_coeff_mult_21_n106), .ZN(
        my_filter_first_coeff_mult_21_ab_7__9_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U101 ( .A1(
        my_filter_first_coeff_mult_21_n92), .A2(
        my_filter_first_coeff_mult_21_n106), .ZN(
        my_filter_first_coeff_mult_21_ab_7__7_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U100 ( .A1(
        my_filter_first_coeff_mult_21_n97), .A2(
        my_filter_first_coeff_mult_21_n105), .ZN(
        my_filter_first_coeff_mult_21_ab_8__2_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U99 ( .A1(
        my_filter_first_coeff_mult_21_n95), .A2(
        my_filter_first_coeff_mult_21_n105), .ZN(
        my_filter_first_coeff_mult_21_ab_8__4_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U98 ( .A1(
        my_filter_first_coeff_mult_21_n94), .A2(
        my_filter_first_coeff_mult_21_n105), .ZN(
        my_filter_first_coeff_mult_21_ab_8__5_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U97 ( .A1(
        my_filter_first_coeff_mult_21_n90), .A2(
        my_filter_first_coeff_mult_21_n107), .ZN(
        my_filter_first_coeff_mult_21_ab_6__9_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U96 ( .A1(
        my_filter_first_coeff_mult_21_n89), .A2(
        my_filter_first_coeff_mult_21_n107), .ZN(
        my_filter_first_coeff_mult_21_ab_6__10_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U95 ( .A1(
        my_filter_first_coeff_mult_21_n91), .A2(
        my_filter_first_coeff_mult_21_n107), .ZN(
        my_filter_first_coeff_mult_21_ab_6__8_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U94 ( .A1(
        my_filter_first_coeff_mult_21_n93), .A2(
        my_filter_first_coeff_mult_21_n106), .ZN(
        my_filter_first_coeff_mult_21_ab_7__6_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U93 ( .A1(
        my_filter_first_coeff_mult_21_n89), .A2(
        my_filter_first_coeff_mult_21_n108), .ZN(
        my_filter_first_coeff_mult_21_ab_5__10_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U92 ( .A1(
        my_filter_first_coeff_mult_21_n88), .A2(
        my_filter_first_coeff_mult_21_n108), .ZN(
        my_filter_first_coeff_mult_21_ab_5__11_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U91 ( .A1(
        my_filter_first_coeff_mult_21_n90), .A2(
        my_filter_first_coeff_mult_21_n108), .ZN(
        my_filter_first_coeff_mult_21_ab_5__9_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U90 ( .A1(
        my_filter_first_coeff_mult_21_n97), .A2(
        my_filter_first_coeff_mult_21_n107), .ZN(
        my_filter_first_coeff_mult_21_ab_6__2_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U89 ( .A1(
        my_filter_first_coeff_mult_21_n95), .A2(
        my_filter_first_coeff_mult_21_n107), .ZN(
        my_filter_first_coeff_mult_21_ab_6__4_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U88 ( .A1(
        my_filter_first_coeff_mult_21_n93), .A2(
        my_filter_first_coeff_mult_21_n107), .ZN(
        my_filter_first_coeff_mult_21_ab_6__6_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U87 ( .A1(
        my_filter_first_coeff_mult_21_n92), .A2(
        my_filter_first_coeff_mult_21_n107), .ZN(
        my_filter_first_coeff_mult_21_ab_6__7_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U86 ( .A1(
        my_filter_first_coeff_mult_21_n88), .A2(
        my_filter_first_coeff_mult_21_n109), .ZN(
        my_filter_first_coeff_mult_21_ab_4__11_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U85 ( .A1(
        my_filter_first_coeff_mult_21_n89), .A2(
        my_filter_first_coeff_mult_21_n109), .ZN(
        my_filter_first_coeff_mult_21_ab_4__10_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U84 ( .A1(
        my_filter_first_coeff_mult_21_n91), .A2(
        my_filter_first_coeff_mult_21_n108), .ZN(
        my_filter_first_coeff_mult_21_ab_5__8_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U83 ( .A1(
        my_filter_first_coeff_mult_21_n88), .A2(
        my_filter_first_coeff_mult_21_n110), .ZN(
        my_filter_first_coeff_mult_21_ab_3__11_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U82 ( .A1(
        my_filter_first_coeff_mult_21_n97), .A2(
        my_filter_first_coeff_mult_21_n109), .ZN(
        my_filter_first_coeff_mult_21_ab_4__2_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U81 ( .A1(
        my_filter_first_coeff_mult_21_n95), .A2(
        my_filter_first_coeff_mult_21_n109), .ZN(
        my_filter_first_coeff_mult_21_ab_4__4_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U80 ( .A1(
        my_filter_first_coeff_mult_21_n93), .A2(
        my_filter_first_coeff_mult_21_n109), .ZN(
        my_filter_first_coeff_mult_21_ab_4__6_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U79 ( .A1(
        my_filter_first_coeff_mult_21_n92), .A2(
        my_filter_first_coeff_mult_21_n109), .ZN(
        my_filter_first_coeff_mult_21_ab_4__7_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U78 ( .A1(
        my_filter_first_coeff_mult_21_n91), .A2(
        my_filter_first_coeff_mult_21_n109), .ZN(
        my_filter_first_coeff_mult_21_ab_4__8_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U77 ( .A1(
        my_filter_first_coeff_mult_21_n90), .A2(
        my_filter_first_coeff_mult_21_n109), .ZN(
        my_filter_first_coeff_mult_21_ab_4__9_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U76 ( .A1(
        my_filter_first_coeff_mult_21_n92), .A2(
        my_filter_first_coeff_mult_21_n110), .ZN(
        my_filter_first_coeff_mult_21_ab_3__7_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U75 ( .A1(
        my_filter_first_coeff_mult_21_n89), .A2(
        my_filter_first_coeff_mult_21_n110), .ZN(
        my_filter_first_coeff_mult_21_ab_3__10_) );
  AND2_X1 my_filter_first_coeff_mult_21_U74 ( .A1(
        my_filter_first_coeff_mult_21_ab_0__2_), .A2(
        my_filter_first_coeff_mult_21_ab_1__1_), .ZN(
        my_filter_first_coeff_mult_21_n14) );
  NOR2_X1 my_filter_first_coeff_mult_21_U73 ( .A1(
        my_filter_first_coeff_mult_21_n98), .A2(
        my_filter_first_coeff_mult_21_n111), .ZN(
        my_filter_first_coeff_mult_21_ab_2__1_) );
  AND2_X1 my_filter_first_coeff_mult_21_U72 ( .A1(
        my_filter_first_coeff_mult_21_ab_0__3_), .A2(
        my_filter_first_coeff_mult_21_ab_1__2_), .ZN(
        my_filter_first_coeff_mult_21_n13) );
  NOR2_X1 my_filter_first_coeff_mult_21_U71 ( .A1(
        my_filter_first_coeff_mult_21_n97), .A2(
        my_filter_first_coeff_mult_21_n111), .ZN(
        my_filter_first_coeff_mult_21_ab_2__2_) );
  AND2_X1 my_filter_first_coeff_mult_21_U70 ( .A1(
        my_filter_first_coeff_mult_21_ab_0__4_), .A2(
        my_filter_first_coeff_mult_21_ab_1__3_), .ZN(
        my_filter_first_coeff_mult_21_n12) );
  NOR2_X1 my_filter_first_coeff_mult_21_U69 ( .A1(
        my_filter_first_coeff_mult_21_n96), .A2(
        my_filter_first_coeff_mult_21_n111), .ZN(
        my_filter_first_coeff_mult_21_ab_2__3_) );
  AND2_X1 my_filter_first_coeff_mult_21_U68 ( .A1(
        my_filter_first_coeff_mult_21_ab_0__5_), .A2(
        my_filter_first_coeff_mult_21_ab_1__4_), .ZN(
        my_filter_first_coeff_mult_21_n11) );
  NOR2_X1 my_filter_first_coeff_mult_21_U67 ( .A1(
        my_filter_first_coeff_mult_21_n95), .A2(
        my_filter_first_coeff_mult_21_n111), .ZN(
        my_filter_first_coeff_mult_21_ab_2__4_) );
  AND2_X1 my_filter_first_coeff_mult_21_U66 ( .A1(
        my_filter_first_coeff_mult_21_ab_0__6_), .A2(
        my_filter_first_coeff_mult_21_ab_1__5_), .ZN(
        my_filter_first_coeff_mult_21_n10) );
  NOR2_X1 my_filter_first_coeff_mult_21_U65 ( .A1(
        my_filter_first_coeff_mult_21_n94), .A2(
        my_filter_first_coeff_mult_21_n111), .ZN(
        my_filter_first_coeff_mult_21_ab_2__5_) );
  AND2_X1 my_filter_first_coeff_mult_21_U64 ( .A1(
        my_filter_first_coeff_mult_21_ab_0__7_), .A2(
        my_filter_first_coeff_mult_21_ab_1__6_), .ZN(
        my_filter_first_coeff_mult_21_n9) );
  NOR2_X1 my_filter_first_coeff_mult_21_U63 ( .A1(
        my_filter_first_coeff_mult_21_n93), .A2(
        my_filter_first_coeff_mult_21_n111), .ZN(
        my_filter_first_coeff_mult_21_ab_2__6_) );
  AND2_X1 my_filter_first_coeff_mult_21_U62 ( .A1(
        my_filter_first_coeff_mult_21_ab_0__8_), .A2(
        my_filter_first_coeff_mult_21_ab_1__7_), .ZN(
        my_filter_first_coeff_mult_21_n8) );
  NOR2_X1 my_filter_first_coeff_mult_21_U61 ( .A1(
        my_filter_first_coeff_mult_21_n92), .A2(
        my_filter_first_coeff_mult_21_n111), .ZN(
        my_filter_first_coeff_mult_21_ab_2__7_) );
  AND2_X1 my_filter_first_coeff_mult_21_U60 ( .A1(
        my_filter_first_coeff_mult_21_ab_0__9_), .A2(
        my_filter_first_coeff_mult_21_ab_1__8_), .ZN(
        my_filter_first_coeff_mult_21_n7) );
  NOR2_X1 my_filter_first_coeff_mult_21_U59 ( .A1(
        my_filter_first_coeff_mult_21_n91), .A2(
        my_filter_first_coeff_mult_21_n111), .ZN(
        my_filter_first_coeff_mult_21_ab_2__8_) );
  AND2_X1 my_filter_first_coeff_mult_21_U58 ( .A1(
        my_filter_first_coeff_mult_21_ab_0__10_), .A2(
        my_filter_first_coeff_mult_21_ab_1__9_), .ZN(
        my_filter_first_coeff_mult_21_n6) );
  NOR2_X1 my_filter_first_coeff_mult_21_U57 ( .A1(
        my_filter_first_coeff_mult_21_n90), .A2(
        my_filter_first_coeff_mult_21_n111), .ZN(
        my_filter_first_coeff_mult_21_ab_2__9_) );
  AND2_X1 my_filter_first_coeff_mult_21_U56 ( .A1(
        my_filter_first_coeff_mult_21_ab_0__11_), .A2(
        my_filter_first_coeff_mult_21_ab_1__10_), .ZN(
        my_filter_first_coeff_mult_21_n5) );
  NOR2_X1 my_filter_first_coeff_mult_21_U55 ( .A1(
        my_filter_first_coeff_mult_21_n89), .A2(
        my_filter_first_coeff_mult_21_n111), .ZN(
        my_filter_first_coeff_mult_21_ab_2__10_) );
  AND2_X1 my_filter_first_coeff_mult_21_U54 ( .A1(
        my_filter_first_coeff_mult_21_ab_0__12_), .A2(
        my_filter_first_coeff_mult_21_ab_1__11_), .ZN(
        my_filter_first_coeff_mult_21_n4) );
  NOR2_X1 my_filter_first_coeff_mult_21_U52 ( .A1(
        my_filter_first_coeff_mult_21_n88), .A2(
        my_filter_first_coeff_mult_21_n111), .ZN(
        my_filter_first_coeff_mult_21_ab_2__11_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U51 ( .A1(
        my_filter_first_coeff_mult_21_n87), .A2(
        my_filter_first_coeff_mult_21_n112), .ZN(
        my_filter_first_coeff_mult_21_ab_1__12_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U49 ( .A1(
        my_filter_first_coeff_mult_21_n97), .A2(
        my_filter_first_coeff_mult_21_n112), .ZN(
        my_filter_first_coeff_mult_21_ab_1__2_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U48 ( .A1(
        my_filter_first_coeff_mult_21_n96), .A2(
        my_filter_first_coeff_mult_21_n112), .ZN(
        my_filter_first_coeff_mult_21_ab_1__3_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U43 ( .A1(
        my_filter_first_coeff_mult_21_n95), .A2(
        my_filter_first_coeff_mult_21_n112), .ZN(
        my_filter_first_coeff_mult_21_ab_1__4_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U42 ( .A1(
        my_filter_first_coeff_mult_21_n94), .A2(
        my_filter_first_coeff_mult_21_n112), .ZN(
        my_filter_first_coeff_mult_21_ab_1__5_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U41 ( .A1(
        my_filter_first_coeff_mult_21_n93), .A2(
        my_filter_first_coeff_mult_21_n112), .ZN(
        my_filter_first_coeff_mult_21_ab_1__6_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U40 ( .A1(
        my_filter_first_coeff_mult_21_n92), .A2(
        my_filter_first_coeff_mult_21_n112), .ZN(
        my_filter_first_coeff_mult_21_ab_1__7_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U39 ( .A1(
        my_filter_first_coeff_mult_21_n91), .A2(
        my_filter_first_coeff_mult_21_n112), .ZN(
        my_filter_first_coeff_mult_21_ab_1__8_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U38 ( .A1(
        my_filter_first_coeff_mult_21_n90), .A2(
        my_filter_first_coeff_mult_21_n112), .ZN(
        my_filter_first_coeff_mult_21_ab_1__9_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U34 ( .A1(
        my_filter_first_coeff_mult_21_n89), .A2(
        my_filter_first_coeff_mult_21_n112), .ZN(
        my_filter_first_coeff_mult_21_ab_1__10_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U26 ( .A1(
        my_filter_first_coeff_mult_21_n88), .A2(
        my_filter_first_coeff_mult_21_n112), .ZN(
        my_filter_first_coeff_mult_21_ab_1__11_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U14 ( .A1(
        my_filter_first_coeff_mult_21_n97), .A2(
        my_filter_first_coeff_mult_21_n113), .ZN(
        my_filter_first_coeff_mult_21_ab_0__2_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U13 ( .A1(
        my_filter_first_coeff_mult_21_n96), .A2(
        my_filter_first_coeff_mult_21_n113), .ZN(
        my_filter_first_coeff_mult_21_ab_0__3_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U12 ( .A1(
        my_filter_first_coeff_mult_21_n95), .A2(
        my_filter_first_coeff_mult_21_n113), .ZN(
        my_filter_first_coeff_mult_21_ab_0__4_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U11 ( .A1(
        my_filter_first_coeff_mult_21_n94), .A2(
        my_filter_first_coeff_mult_21_n113), .ZN(
        my_filter_first_coeff_mult_21_ab_0__5_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U10 ( .A1(
        my_filter_first_coeff_mult_21_n93), .A2(
        my_filter_first_coeff_mult_21_n113), .ZN(
        my_filter_first_coeff_mult_21_ab_0__6_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U9 ( .A1(
        my_filter_first_coeff_mult_21_n92), .A2(
        my_filter_first_coeff_mult_21_n113), .ZN(
        my_filter_first_coeff_mult_21_ab_0__7_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U8 ( .A1(
        my_filter_first_coeff_mult_21_n91), .A2(
        my_filter_first_coeff_mult_21_n113), .ZN(
        my_filter_first_coeff_mult_21_ab_0__8_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U7 ( .A1(
        my_filter_first_coeff_mult_21_n90), .A2(
        my_filter_first_coeff_mult_21_n113), .ZN(
        my_filter_first_coeff_mult_21_ab_0__9_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U6 ( .A1(
        my_filter_first_coeff_mult_21_n89), .A2(
        my_filter_first_coeff_mult_21_n113), .ZN(
        my_filter_first_coeff_mult_21_ab_0__10_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U5 ( .A1(
        my_filter_first_coeff_mult_21_n88), .A2(
        my_filter_first_coeff_mult_21_n113), .ZN(
        my_filter_first_coeff_mult_21_ab_0__11_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U4 ( .A1(
        my_filter_first_coeff_mult_21_n87), .A2(
        my_filter_first_coeff_mult_21_n113), .ZN(
        my_filter_first_coeff_mult_21_ab_0__12_) );
  NOR2_X1 my_filter_first_coeff_mult_21_U3 ( .A1(
        my_filter_first_coeff_mult_21_n112), .A2(
        my_filter_first_coeff_mult_21_n98), .ZN(
        my_filter_first_coeff_mult_21_ab_1__1_) );
  INV_X1 my_filter_first_coeff_mult_21_U2 ( .A(
        my_filter_first_coeff_mult_21_CARRYB_13__13_), .ZN(
        my_filter_first_coeff_mult_21_n85) );
  XOR2_X1 my_filter_first_coeff_mult_21_U50 ( .A(
        my_filter_first_coeff_mult_21_CARRYB_13__10_), .B(
        my_filter_first_coeff_mult_21_SUMB_13__11_), .Z(
        my_filter_first_coeff_mult_21_n50) );
  XOR2_X1 my_filter_first_coeff_mult_21_U47 ( .A(
        my_filter_first_coeff_mult_21_CARRYB_13__11_), .B(
        my_filter_first_coeff_mult_21_SUMB_13__12_), .Z(
        my_filter_first_coeff_mult_21_n47) );
  XOR2_X1 my_filter_first_coeff_mult_21_U46 ( .A(
        my_filter_first_coeff_mult_21_CARRYB_13__8_), .B(
        my_filter_first_coeff_mult_21_SUMB_13__9_), .Z(
        my_filter_first_coeff_mult_21_n46) );
  XOR2_X1 my_filter_first_coeff_mult_21_U45 ( .A(
        my_filter_first_coeff_mult_21_CARRYB_13__9_), .B(
        my_filter_first_coeff_mult_21_SUMB_13__10_), .Z(
        my_filter_first_coeff_mult_21_n45) );
  XOR2_X1 my_filter_first_coeff_mult_21_U44 ( .A(
        my_filter_first_coeff_mult_21_CARRYB_13__12_), .B(
        my_filter_first_coeff_mult_21_SUMB_13__13_), .Z(
        my_filter_first_coeff_mult_21_n44) );
  XOR2_X1 my_filter_first_coeff_mult_21_U37 ( .A(
        my_filter_first_coeff_mult_21_CARRYB_13__5_), .B(
        my_filter_first_coeff_mult_21_SUMB_13__6_), .Z(
        my_filter_first_coeff_mult_21_n37) );
  XOR2_X1 my_filter_first_coeff_mult_21_U36 ( .A(
        my_filter_first_coeff_mult_21_CARRYB_13__3_), .B(
        my_filter_first_coeff_mult_21_SUMB_13__4_), .Z(
        my_filter_first_coeff_mult_21_n36) );
  XOR2_X1 my_filter_first_coeff_mult_21_U35 ( .A(
        my_filter_first_coeff_mult_21_CARRYB_13__1_), .B(
        my_filter_first_coeff_mult_21_SUMB_13__2_), .Z(
        my_filter_first_coeff_mult_21_n35) );
  XOR2_X1 my_filter_first_coeff_mult_21_U33 ( .A(
        my_filter_first_coeff_mult_21_CARRYB_13__6_), .B(
        my_filter_first_coeff_mult_21_SUMB_13__7_), .Z(
        my_filter_first_coeff_mult_21_n33) );
  XOR2_X1 my_filter_first_coeff_mult_21_U32 ( .A(
        my_filter_first_coeff_mult_21_CARRYB_13__7_), .B(
        my_filter_first_coeff_mult_21_SUMB_13__8_), .Z(
        my_filter_first_coeff_mult_21_n32) );
  XOR2_X1 my_filter_first_coeff_mult_21_U31 ( .A(
        my_filter_first_coeff_mult_21_CARRYB_13__4_), .B(
        my_filter_first_coeff_mult_21_SUMB_13__5_), .Z(
        my_filter_first_coeff_mult_21_n31) );
  XOR2_X1 my_filter_first_coeff_mult_21_U30 ( .A(
        my_filter_first_coeff_mult_21_CARRYB_13__2_), .B(
        my_filter_first_coeff_mult_21_SUMB_13__3_), .Z(
        my_filter_first_coeff_mult_21_n30) );
  XOR2_X1 my_filter_first_coeff_mult_21_U29 ( .A(
        my_filter_first_coeff_mult_21_CARRYB_13__0_), .B(
        my_filter_first_coeff_mult_21_SUMB_13__1_), .Z(
        my_filter_first_coeff_mult_21_n29) );
  XOR2_X1 my_filter_first_coeff_mult_21_U27 ( .A(
        my_filter_first_coeff_mult_21_ab_1__1_), .B(
        my_filter_first_coeff_mult_21_ab_0__2_), .Z(
        my_filter_first_coeff_mult_21_n28) );
  XOR2_X1 my_filter_first_coeff_mult_21_U25 ( .A(
        my_filter_first_coeff_mult_21_ab_1__12_), .B(
        my_filter_first_coeff_mult_21_ab_0__13_), .Z(
        my_filter_first_coeff_mult_21_n26) );
  XOR2_X1 my_filter_first_coeff_mult_21_U24 ( .A(
        my_filter_first_coeff_mult_21_ab_1__2_), .B(
        my_filter_first_coeff_mult_21_ab_0__3_), .Z(
        my_filter_first_coeff_mult_21_n25) );
  XOR2_X1 my_filter_first_coeff_mult_21_U23 ( .A(
        my_filter_first_coeff_mult_21_ab_1__3_), .B(
        my_filter_first_coeff_mult_21_ab_0__4_), .Z(
        my_filter_first_coeff_mult_21_n24) );
  XOR2_X1 my_filter_first_coeff_mult_21_U22 ( .A(
        my_filter_first_coeff_mult_21_ab_1__4_), .B(
        my_filter_first_coeff_mult_21_ab_0__5_), .Z(
        my_filter_first_coeff_mult_21_n23) );
  XOR2_X1 my_filter_first_coeff_mult_21_U21 ( .A(
        my_filter_first_coeff_mult_21_ab_1__5_), .B(
        my_filter_first_coeff_mult_21_ab_0__6_), .Z(
        my_filter_first_coeff_mult_21_n22) );
  XOR2_X1 my_filter_first_coeff_mult_21_U20 ( .A(
        my_filter_first_coeff_mult_21_ab_1__6_), .B(
        my_filter_first_coeff_mult_21_ab_0__7_), .Z(
        my_filter_first_coeff_mult_21_n21) );
  XOR2_X1 my_filter_first_coeff_mult_21_U19 ( .A(
        my_filter_first_coeff_mult_21_ab_1__7_), .B(
        my_filter_first_coeff_mult_21_ab_0__8_), .Z(
        my_filter_first_coeff_mult_21_n20) );
  XOR2_X1 my_filter_first_coeff_mult_21_U18 ( .A(
        my_filter_first_coeff_mult_21_ab_1__8_), .B(
        my_filter_first_coeff_mult_21_ab_0__9_), .Z(
        my_filter_first_coeff_mult_21_n19) );
  XOR2_X1 my_filter_first_coeff_mult_21_U17 ( .A(
        my_filter_first_coeff_mult_21_ab_1__9_), .B(
        my_filter_first_coeff_mult_21_ab_0__10_), .Z(
        my_filter_first_coeff_mult_21_n18) );
  XOR2_X1 my_filter_first_coeff_mult_21_U16 ( .A(
        my_filter_first_coeff_mult_21_ab_1__10_), .B(
        my_filter_first_coeff_mult_21_ab_0__11_), .Z(
        my_filter_first_coeff_mult_21_n17) );
  XOR2_X1 my_filter_first_coeff_mult_21_U15 ( .A(
        my_filter_first_coeff_mult_21_ab_1__11_), .B(
        my_filter_first_coeff_mult_21_ab_0__12_), .Z(
        my_filter_first_coeff_mult_21_n16) );
  FA_X1 my_filter_first_coeff_mult_21_S3_2_12 ( .A(
        my_filter_first_coeff_mult_21_ab_2__12_), .B(
        my_filter_first_coeff_mult_21_n15), .CI(
        my_filter_first_coeff_mult_21_ab_1__13_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_2__12_), .S(
        my_filter_first_coeff_mult_21_SUMB_2__12_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_2_11 ( .A(
        my_filter_first_coeff_mult_21_ab_2__11_), .B(
        my_filter_first_coeff_mult_21_n4), .CI(
        my_filter_first_coeff_mult_21_n26), .CO(
        my_filter_first_coeff_mult_21_CARRYB_2__11_), .S(
        my_filter_first_coeff_mult_21_SUMB_2__11_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_2_10 ( .A(
        my_filter_first_coeff_mult_21_ab_2__10_), .B(
        my_filter_first_coeff_mult_21_n5), .CI(
        my_filter_first_coeff_mult_21_n16), .CO(
        my_filter_first_coeff_mult_21_CARRYB_2__10_), .S(
        my_filter_first_coeff_mult_21_SUMB_2__10_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_2_9 ( .A(
        my_filter_first_coeff_mult_21_ab_2__9_), .B(
        my_filter_first_coeff_mult_21_n6), .CI(
        my_filter_first_coeff_mult_21_n17), .CO(
        my_filter_first_coeff_mult_21_CARRYB_2__9_), .S(
        my_filter_first_coeff_mult_21_SUMB_2__9_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_2_8 ( .A(
        my_filter_first_coeff_mult_21_ab_2__8_), .B(
        my_filter_first_coeff_mult_21_n7), .CI(
        my_filter_first_coeff_mult_21_n18), .CO(
        my_filter_first_coeff_mult_21_CARRYB_2__8_), .S(
        my_filter_first_coeff_mult_21_SUMB_2__8_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_2_7 ( .A(
        my_filter_first_coeff_mult_21_ab_2__7_), .B(
        my_filter_first_coeff_mult_21_n8), .CI(
        my_filter_first_coeff_mult_21_n19), .CO(
        my_filter_first_coeff_mult_21_CARRYB_2__7_), .S(
        my_filter_first_coeff_mult_21_SUMB_2__7_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_2_6 ( .A(
        my_filter_first_coeff_mult_21_ab_2__6_), .B(
        my_filter_first_coeff_mult_21_n9), .CI(
        my_filter_first_coeff_mult_21_n20), .CO(
        my_filter_first_coeff_mult_21_CARRYB_2__6_), .S(
        my_filter_first_coeff_mult_21_SUMB_2__6_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_2_5 ( .A(
        my_filter_first_coeff_mult_21_ab_2__5_), .B(
        my_filter_first_coeff_mult_21_n10), .CI(
        my_filter_first_coeff_mult_21_n21), .CO(
        my_filter_first_coeff_mult_21_CARRYB_2__5_), .S(
        my_filter_first_coeff_mult_21_SUMB_2__5_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_2_4 ( .A(
        my_filter_first_coeff_mult_21_ab_2__4_), .B(
        my_filter_first_coeff_mult_21_n11), .CI(
        my_filter_first_coeff_mult_21_n22), .CO(
        my_filter_first_coeff_mult_21_CARRYB_2__4_), .S(
        my_filter_first_coeff_mult_21_SUMB_2__4_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_2_3 ( .A(
        my_filter_first_coeff_mult_21_ab_2__3_), .B(
        my_filter_first_coeff_mult_21_n12), .CI(
        my_filter_first_coeff_mult_21_n23), .CO(
        my_filter_first_coeff_mult_21_CARRYB_2__3_), .S(
        my_filter_first_coeff_mult_21_SUMB_2__3_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_2_2 ( .A(
        my_filter_first_coeff_mult_21_ab_2__2_), .B(
        my_filter_first_coeff_mult_21_n13), .CI(
        my_filter_first_coeff_mult_21_n24), .CO(
        my_filter_first_coeff_mult_21_CARRYB_2__2_), .S(
        my_filter_first_coeff_mult_21_SUMB_2__2_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_2_1 ( .A(
        my_filter_first_coeff_mult_21_ab_2__1_), .B(
        my_filter_first_coeff_mult_21_n14), .CI(
        my_filter_first_coeff_mult_21_n25), .CO(
        my_filter_first_coeff_mult_21_CARRYB_2__1_), .S(
        my_filter_first_coeff_mult_21_SUMB_2__1_) );
  FA_X1 my_filter_first_coeff_mult_21_S1_2_0 ( .A(
        my_filter_first_coeff_mult_21_ab_2__0_), .B(
        my_filter_first_coeff_mult_21_CARRYB_1__0_), .CI(
        my_filter_first_coeff_mult_21_n28), .CO(
        my_filter_first_coeff_mult_21_CARRYB_2__0_), .S(
        my_filter_first_coeff_mult_21_A1_0_) );
  FA_X1 my_filter_first_coeff_mult_21_S3_3_12 ( .A(
        my_filter_first_coeff_mult_21_ab_3__12_), .B(
        my_filter_first_coeff_mult_21_CARRYB_2__12_), .CI(
        my_filter_first_coeff_mult_21_ab_2__13_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_3__12_), .S(
        my_filter_first_coeff_mult_21_SUMB_3__12_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_3_11 ( .A(
        my_filter_first_coeff_mult_21_ab_3__11_), .B(
        my_filter_first_coeff_mult_21_CARRYB_2__11_), .CI(
        my_filter_first_coeff_mult_21_SUMB_2__12_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_3__11_), .S(
        my_filter_first_coeff_mult_21_SUMB_3__11_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_3_10 ( .A(
        my_filter_first_coeff_mult_21_ab_3__10_), .B(
        my_filter_first_coeff_mult_21_CARRYB_2__10_), .CI(
        my_filter_first_coeff_mult_21_SUMB_2__11_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_3__10_), .S(
        my_filter_first_coeff_mult_21_SUMB_3__10_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_3_9 ( .A(
        my_filter_first_coeff_mult_21_ab_3__9_), .B(
        my_filter_first_coeff_mult_21_CARRYB_2__9_), .CI(
        my_filter_first_coeff_mult_21_SUMB_2__10_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_3__9_), .S(
        my_filter_first_coeff_mult_21_SUMB_3__9_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_3_8 ( .A(
        my_filter_first_coeff_mult_21_ab_3__8_), .B(
        my_filter_first_coeff_mult_21_CARRYB_2__8_), .CI(
        my_filter_first_coeff_mult_21_SUMB_2__9_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_3__8_), .S(
        my_filter_first_coeff_mult_21_SUMB_3__8_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_3_7 ( .A(
        my_filter_first_coeff_mult_21_ab_3__7_), .B(
        my_filter_first_coeff_mult_21_CARRYB_2__7_), .CI(
        my_filter_first_coeff_mult_21_SUMB_2__8_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_3__7_), .S(
        my_filter_first_coeff_mult_21_SUMB_3__7_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_3_6 ( .A(
        my_filter_first_coeff_mult_21_ab_3__6_), .B(
        my_filter_first_coeff_mult_21_CARRYB_2__6_), .CI(
        my_filter_first_coeff_mult_21_SUMB_2__7_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_3__6_), .S(
        my_filter_first_coeff_mult_21_SUMB_3__6_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_3_5 ( .A(
        my_filter_first_coeff_mult_21_ab_3__5_), .B(
        my_filter_first_coeff_mult_21_CARRYB_2__5_), .CI(
        my_filter_first_coeff_mult_21_SUMB_2__6_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_3__5_), .S(
        my_filter_first_coeff_mult_21_SUMB_3__5_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_3_4 ( .A(
        my_filter_first_coeff_mult_21_ab_3__4_), .B(
        my_filter_first_coeff_mult_21_CARRYB_2__4_), .CI(
        my_filter_first_coeff_mult_21_SUMB_2__5_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_3__4_), .S(
        my_filter_first_coeff_mult_21_SUMB_3__4_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_3_3 ( .A(
        my_filter_first_coeff_mult_21_ab_3__3_), .B(
        my_filter_first_coeff_mult_21_CARRYB_2__3_), .CI(
        my_filter_first_coeff_mult_21_SUMB_2__4_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_3__3_), .S(
        my_filter_first_coeff_mult_21_SUMB_3__3_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_3_2 ( .A(
        my_filter_first_coeff_mult_21_ab_3__2_), .B(
        my_filter_first_coeff_mult_21_CARRYB_2__2_), .CI(
        my_filter_first_coeff_mult_21_SUMB_2__3_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_3__2_), .S(
        my_filter_first_coeff_mult_21_SUMB_3__2_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_3_1 ( .A(
        my_filter_first_coeff_mult_21_ab_3__1_), .B(
        my_filter_first_coeff_mult_21_CARRYB_2__1_), .CI(
        my_filter_first_coeff_mult_21_SUMB_2__2_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_3__1_), .S(
        my_filter_first_coeff_mult_21_SUMB_3__1_) );
  FA_X1 my_filter_first_coeff_mult_21_S1_3_0 ( .A(
        my_filter_first_coeff_mult_21_ab_3__0_), .B(
        my_filter_first_coeff_mult_21_CARRYB_2__0_), .CI(
        my_filter_first_coeff_mult_21_SUMB_2__1_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_3__0_), .S(
        my_filter_first_coeff_mult_21_A1_1_) );
  FA_X1 my_filter_first_coeff_mult_21_S3_4_12 ( .A(
        my_filter_first_coeff_mult_21_ab_4__12_), .B(
        my_filter_first_coeff_mult_21_CARRYB_3__12_), .CI(
        my_filter_first_coeff_mult_21_ab_3__13_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_4__12_), .S(
        my_filter_first_coeff_mult_21_SUMB_4__12_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_4_11 ( .A(
        my_filter_first_coeff_mult_21_ab_4__11_), .B(
        my_filter_first_coeff_mult_21_CARRYB_3__11_), .CI(
        my_filter_first_coeff_mult_21_SUMB_3__12_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_4__11_), .S(
        my_filter_first_coeff_mult_21_SUMB_4__11_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_4_10 ( .A(
        my_filter_first_coeff_mult_21_ab_4__10_), .B(
        my_filter_first_coeff_mult_21_CARRYB_3__10_), .CI(
        my_filter_first_coeff_mult_21_SUMB_3__11_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_4__10_), .S(
        my_filter_first_coeff_mult_21_SUMB_4__10_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_4_9 ( .A(
        my_filter_first_coeff_mult_21_ab_4__9_), .B(
        my_filter_first_coeff_mult_21_CARRYB_3__9_), .CI(
        my_filter_first_coeff_mult_21_SUMB_3__10_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_4__9_), .S(
        my_filter_first_coeff_mult_21_SUMB_4__9_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_4_8 ( .A(
        my_filter_first_coeff_mult_21_ab_4__8_), .B(
        my_filter_first_coeff_mult_21_CARRYB_3__8_), .CI(
        my_filter_first_coeff_mult_21_SUMB_3__9_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_4__8_), .S(
        my_filter_first_coeff_mult_21_SUMB_4__8_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_4_7 ( .A(
        my_filter_first_coeff_mult_21_ab_4__7_), .B(
        my_filter_first_coeff_mult_21_CARRYB_3__7_), .CI(
        my_filter_first_coeff_mult_21_SUMB_3__8_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_4__7_), .S(
        my_filter_first_coeff_mult_21_SUMB_4__7_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_4_6 ( .A(
        my_filter_first_coeff_mult_21_ab_4__6_), .B(
        my_filter_first_coeff_mult_21_CARRYB_3__6_), .CI(
        my_filter_first_coeff_mult_21_SUMB_3__7_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_4__6_), .S(
        my_filter_first_coeff_mult_21_SUMB_4__6_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_4_5 ( .A(
        my_filter_first_coeff_mult_21_ab_4__5_), .B(
        my_filter_first_coeff_mult_21_CARRYB_3__5_), .CI(
        my_filter_first_coeff_mult_21_SUMB_3__6_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_4__5_), .S(
        my_filter_first_coeff_mult_21_SUMB_4__5_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_4_4 ( .A(
        my_filter_first_coeff_mult_21_ab_4__4_), .B(
        my_filter_first_coeff_mult_21_CARRYB_3__4_), .CI(
        my_filter_first_coeff_mult_21_SUMB_3__5_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_4__4_), .S(
        my_filter_first_coeff_mult_21_SUMB_4__4_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_4_3 ( .A(
        my_filter_first_coeff_mult_21_ab_4__3_), .B(
        my_filter_first_coeff_mult_21_CARRYB_3__3_), .CI(
        my_filter_first_coeff_mult_21_SUMB_3__4_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_4__3_), .S(
        my_filter_first_coeff_mult_21_SUMB_4__3_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_4_2 ( .A(
        my_filter_first_coeff_mult_21_ab_4__2_), .B(
        my_filter_first_coeff_mult_21_CARRYB_3__2_), .CI(
        my_filter_first_coeff_mult_21_SUMB_3__3_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_4__2_), .S(
        my_filter_first_coeff_mult_21_SUMB_4__2_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_4_1 ( .A(
        my_filter_first_coeff_mult_21_ab_4__1_), .B(
        my_filter_first_coeff_mult_21_CARRYB_3__1_), .CI(
        my_filter_first_coeff_mult_21_SUMB_3__2_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_4__1_), .S(
        my_filter_first_coeff_mult_21_SUMB_4__1_) );
  FA_X1 my_filter_first_coeff_mult_21_S1_4_0 ( .A(
        my_filter_first_coeff_mult_21_ab_4__0_), .B(
        my_filter_first_coeff_mult_21_CARRYB_3__0_), .CI(
        my_filter_first_coeff_mult_21_SUMB_3__1_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_4__0_), .S(
        my_filter_first_coeff_mult_21_A1_2_) );
  FA_X1 my_filter_first_coeff_mult_21_S3_5_12 ( .A(
        my_filter_first_coeff_mult_21_ab_5__12_), .B(
        my_filter_first_coeff_mult_21_CARRYB_4__12_), .CI(
        my_filter_first_coeff_mult_21_ab_4__13_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_5__12_), .S(
        my_filter_first_coeff_mult_21_SUMB_5__12_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_5_11 ( .A(
        my_filter_first_coeff_mult_21_ab_5__11_), .B(
        my_filter_first_coeff_mult_21_CARRYB_4__11_), .CI(
        my_filter_first_coeff_mult_21_SUMB_4__12_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_5__11_), .S(
        my_filter_first_coeff_mult_21_SUMB_5__11_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_5_10 ( .A(
        my_filter_first_coeff_mult_21_ab_5__10_), .B(
        my_filter_first_coeff_mult_21_CARRYB_4__10_), .CI(
        my_filter_first_coeff_mult_21_SUMB_4__11_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_5__10_), .S(
        my_filter_first_coeff_mult_21_SUMB_5__10_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_5_9 ( .A(
        my_filter_first_coeff_mult_21_ab_5__9_), .B(
        my_filter_first_coeff_mult_21_CARRYB_4__9_), .CI(
        my_filter_first_coeff_mult_21_SUMB_4__10_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_5__9_), .S(
        my_filter_first_coeff_mult_21_SUMB_5__9_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_5_8 ( .A(
        my_filter_first_coeff_mult_21_ab_5__8_), .B(
        my_filter_first_coeff_mult_21_CARRYB_4__8_), .CI(
        my_filter_first_coeff_mult_21_SUMB_4__9_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_5__8_), .S(
        my_filter_first_coeff_mult_21_SUMB_5__8_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_5_7 ( .A(
        my_filter_first_coeff_mult_21_ab_5__7_), .B(
        my_filter_first_coeff_mult_21_CARRYB_4__7_), .CI(
        my_filter_first_coeff_mult_21_SUMB_4__8_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_5__7_), .S(
        my_filter_first_coeff_mult_21_SUMB_5__7_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_5_6 ( .A(
        my_filter_first_coeff_mult_21_ab_5__6_), .B(
        my_filter_first_coeff_mult_21_CARRYB_4__6_), .CI(
        my_filter_first_coeff_mult_21_SUMB_4__7_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_5__6_), .S(
        my_filter_first_coeff_mult_21_SUMB_5__6_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_5_5 ( .A(
        my_filter_first_coeff_mult_21_ab_5__5_), .B(
        my_filter_first_coeff_mult_21_CARRYB_4__5_), .CI(
        my_filter_first_coeff_mult_21_SUMB_4__6_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_5__5_), .S(
        my_filter_first_coeff_mult_21_SUMB_5__5_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_5_4 ( .A(
        my_filter_first_coeff_mult_21_ab_5__4_), .B(
        my_filter_first_coeff_mult_21_CARRYB_4__4_), .CI(
        my_filter_first_coeff_mult_21_SUMB_4__5_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_5__4_), .S(
        my_filter_first_coeff_mult_21_SUMB_5__4_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_5_3 ( .A(
        my_filter_first_coeff_mult_21_ab_5__3_), .B(
        my_filter_first_coeff_mult_21_CARRYB_4__3_), .CI(
        my_filter_first_coeff_mult_21_SUMB_4__4_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_5__3_), .S(
        my_filter_first_coeff_mult_21_SUMB_5__3_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_5_2 ( .A(
        my_filter_first_coeff_mult_21_ab_5__2_), .B(
        my_filter_first_coeff_mult_21_CARRYB_4__2_), .CI(
        my_filter_first_coeff_mult_21_SUMB_4__3_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_5__2_), .S(
        my_filter_first_coeff_mult_21_SUMB_5__2_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_5_1 ( .A(
        my_filter_first_coeff_mult_21_ab_5__1_), .B(
        my_filter_first_coeff_mult_21_CARRYB_4__1_), .CI(
        my_filter_first_coeff_mult_21_SUMB_4__2_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_5__1_), .S(
        my_filter_first_coeff_mult_21_SUMB_5__1_) );
  FA_X1 my_filter_first_coeff_mult_21_S1_5_0 ( .A(
        my_filter_first_coeff_mult_21_ab_5__0_), .B(
        my_filter_first_coeff_mult_21_CARRYB_4__0_), .CI(
        my_filter_first_coeff_mult_21_SUMB_4__1_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_5__0_), .S(
        my_filter_first_coeff_mult_21_A1_3_) );
  FA_X1 my_filter_first_coeff_mult_21_S3_6_12 ( .A(
        my_filter_first_coeff_mult_21_ab_6__12_), .B(
        my_filter_first_coeff_mult_21_CARRYB_5__12_), .CI(
        my_filter_first_coeff_mult_21_ab_5__13_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_6__12_), .S(
        my_filter_first_coeff_mult_21_SUMB_6__12_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_6_11 ( .A(
        my_filter_first_coeff_mult_21_ab_6__11_), .B(
        my_filter_first_coeff_mult_21_CARRYB_5__11_), .CI(
        my_filter_first_coeff_mult_21_SUMB_5__12_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_6__11_), .S(
        my_filter_first_coeff_mult_21_SUMB_6__11_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_6_10 ( .A(
        my_filter_first_coeff_mult_21_ab_6__10_), .B(
        my_filter_first_coeff_mult_21_CARRYB_5__10_), .CI(
        my_filter_first_coeff_mult_21_SUMB_5__11_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_6__10_), .S(
        my_filter_first_coeff_mult_21_SUMB_6__10_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_6_9 ( .A(
        my_filter_first_coeff_mult_21_ab_6__9_), .B(
        my_filter_first_coeff_mult_21_CARRYB_5__9_), .CI(
        my_filter_first_coeff_mult_21_SUMB_5__10_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_6__9_), .S(
        my_filter_first_coeff_mult_21_SUMB_6__9_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_6_8 ( .A(
        my_filter_first_coeff_mult_21_ab_6__8_), .B(
        my_filter_first_coeff_mult_21_CARRYB_5__8_), .CI(
        my_filter_first_coeff_mult_21_SUMB_5__9_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_6__8_), .S(
        my_filter_first_coeff_mult_21_SUMB_6__8_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_6_7 ( .A(
        my_filter_first_coeff_mult_21_ab_6__7_), .B(
        my_filter_first_coeff_mult_21_CARRYB_5__7_), .CI(
        my_filter_first_coeff_mult_21_SUMB_5__8_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_6__7_), .S(
        my_filter_first_coeff_mult_21_SUMB_6__7_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_6_6 ( .A(
        my_filter_first_coeff_mult_21_ab_6__6_), .B(
        my_filter_first_coeff_mult_21_CARRYB_5__6_), .CI(
        my_filter_first_coeff_mult_21_SUMB_5__7_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_6__6_), .S(
        my_filter_first_coeff_mult_21_SUMB_6__6_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_6_5 ( .A(
        my_filter_first_coeff_mult_21_ab_6__5_), .B(
        my_filter_first_coeff_mult_21_CARRYB_5__5_), .CI(
        my_filter_first_coeff_mult_21_SUMB_5__6_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_6__5_), .S(
        my_filter_first_coeff_mult_21_SUMB_6__5_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_6_4 ( .A(
        my_filter_first_coeff_mult_21_ab_6__4_), .B(
        my_filter_first_coeff_mult_21_CARRYB_5__4_), .CI(
        my_filter_first_coeff_mult_21_SUMB_5__5_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_6__4_), .S(
        my_filter_first_coeff_mult_21_SUMB_6__4_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_6_3 ( .A(
        my_filter_first_coeff_mult_21_ab_6__3_), .B(
        my_filter_first_coeff_mult_21_CARRYB_5__3_), .CI(
        my_filter_first_coeff_mult_21_SUMB_5__4_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_6__3_), .S(
        my_filter_first_coeff_mult_21_SUMB_6__3_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_6_2 ( .A(
        my_filter_first_coeff_mult_21_ab_6__2_), .B(
        my_filter_first_coeff_mult_21_CARRYB_5__2_), .CI(
        my_filter_first_coeff_mult_21_SUMB_5__3_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_6__2_), .S(
        my_filter_first_coeff_mult_21_SUMB_6__2_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_6_1 ( .A(
        my_filter_first_coeff_mult_21_ab_6__1_), .B(
        my_filter_first_coeff_mult_21_CARRYB_5__1_), .CI(
        my_filter_first_coeff_mult_21_SUMB_5__2_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_6__1_), .S(
        my_filter_first_coeff_mult_21_SUMB_6__1_) );
  FA_X1 my_filter_first_coeff_mult_21_S1_6_0 ( .A(
        my_filter_first_coeff_mult_21_ab_6__0_), .B(
        my_filter_first_coeff_mult_21_CARRYB_5__0_), .CI(
        my_filter_first_coeff_mult_21_SUMB_5__1_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_6__0_), .S(
        my_filter_first_coeff_mult_21_A1_4_) );
  FA_X1 my_filter_first_coeff_mult_21_S3_7_12 ( .A(
        my_filter_first_coeff_mult_21_ab_7__12_), .B(
        my_filter_first_coeff_mult_21_CARRYB_6__12_), .CI(
        my_filter_first_coeff_mult_21_ab_6__13_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_7__12_), .S(
        my_filter_first_coeff_mult_21_SUMB_7__12_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_7_11 ( .A(
        my_filter_first_coeff_mult_21_ab_7__11_), .B(
        my_filter_first_coeff_mult_21_CARRYB_6__11_), .CI(
        my_filter_first_coeff_mult_21_SUMB_6__12_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_7__11_), .S(
        my_filter_first_coeff_mult_21_SUMB_7__11_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_7_10 ( .A(
        my_filter_first_coeff_mult_21_ab_7__10_), .B(
        my_filter_first_coeff_mult_21_CARRYB_6__10_), .CI(
        my_filter_first_coeff_mult_21_SUMB_6__11_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_7__10_), .S(
        my_filter_first_coeff_mult_21_SUMB_7__10_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_7_9 ( .A(
        my_filter_first_coeff_mult_21_ab_7__9_), .B(
        my_filter_first_coeff_mult_21_CARRYB_6__9_), .CI(
        my_filter_first_coeff_mult_21_SUMB_6__10_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_7__9_), .S(
        my_filter_first_coeff_mult_21_SUMB_7__9_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_7_8 ( .A(
        my_filter_first_coeff_mult_21_ab_7__8_), .B(
        my_filter_first_coeff_mult_21_CARRYB_6__8_), .CI(
        my_filter_first_coeff_mult_21_SUMB_6__9_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_7__8_), .S(
        my_filter_first_coeff_mult_21_SUMB_7__8_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_7_7 ( .A(
        my_filter_first_coeff_mult_21_ab_7__7_), .B(
        my_filter_first_coeff_mult_21_CARRYB_6__7_), .CI(
        my_filter_first_coeff_mult_21_SUMB_6__8_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_7__7_), .S(
        my_filter_first_coeff_mult_21_SUMB_7__7_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_7_6 ( .A(
        my_filter_first_coeff_mult_21_ab_7__6_), .B(
        my_filter_first_coeff_mult_21_CARRYB_6__6_), .CI(
        my_filter_first_coeff_mult_21_SUMB_6__7_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_7__6_), .S(
        my_filter_first_coeff_mult_21_SUMB_7__6_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_7_5 ( .A(
        my_filter_first_coeff_mult_21_ab_7__5_), .B(
        my_filter_first_coeff_mult_21_CARRYB_6__5_), .CI(
        my_filter_first_coeff_mult_21_SUMB_6__6_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_7__5_), .S(
        my_filter_first_coeff_mult_21_SUMB_7__5_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_7_4 ( .A(
        my_filter_first_coeff_mult_21_ab_7__4_), .B(
        my_filter_first_coeff_mult_21_CARRYB_6__4_), .CI(
        my_filter_first_coeff_mult_21_SUMB_6__5_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_7__4_), .S(
        my_filter_first_coeff_mult_21_SUMB_7__4_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_7_3 ( .A(
        my_filter_first_coeff_mult_21_ab_7__3_), .B(
        my_filter_first_coeff_mult_21_CARRYB_6__3_), .CI(
        my_filter_first_coeff_mult_21_SUMB_6__4_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_7__3_), .S(
        my_filter_first_coeff_mult_21_SUMB_7__3_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_7_2 ( .A(
        my_filter_first_coeff_mult_21_ab_7__2_), .B(
        my_filter_first_coeff_mult_21_CARRYB_6__2_), .CI(
        my_filter_first_coeff_mult_21_SUMB_6__3_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_7__2_), .S(
        my_filter_first_coeff_mult_21_SUMB_7__2_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_7_1 ( .A(
        my_filter_first_coeff_mult_21_ab_7__1_), .B(
        my_filter_first_coeff_mult_21_CARRYB_6__1_), .CI(
        my_filter_first_coeff_mult_21_SUMB_6__2_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_7__1_), .S(
        my_filter_first_coeff_mult_21_SUMB_7__1_) );
  FA_X1 my_filter_first_coeff_mult_21_S1_7_0 ( .A(
        my_filter_first_coeff_mult_21_ab_7__0_), .B(
        my_filter_first_coeff_mult_21_CARRYB_6__0_), .CI(
        my_filter_first_coeff_mult_21_SUMB_6__1_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_7__0_), .S(
        my_filter_first_coeff_mult_21_A1_5_) );
  FA_X1 my_filter_first_coeff_mult_21_S3_8_12 ( .A(
        my_filter_first_coeff_mult_21_ab_8__12_), .B(
        my_filter_first_coeff_mult_21_CARRYB_7__12_), .CI(
        my_filter_first_coeff_mult_21_ab_7__13_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_8__12_), .S(
        my_filter_first_coeff_mult_21_SUMB_8__12_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_8_11 ( .A(
        my_filter_first_coeff_mult_21_ab_8__11_), .B(
        my_filter_first_coeff_mult_21_CARRYB_7__11_), .CI(
        my_filter_first_coeff_mult_21_SUMB_7__12_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_8__11_), .S(
        my_filter_first_coeff_mult_21_SUMB_8__11_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_8_10 ( .A(
        my_filter_first_coeff_mult_21_ab_8__10_), .B(
        my_filter_first_coeff_mult_21_CARRYB_7__10_), .CI(
        my_filter_first_coeff_mult_21_SUMB_7__11_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_8__10_), .S(
        my_filter_first_coeff_mult_21_SUMB_8__10_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_8_9 ( .A(
        my_filter_first_coeff_mult_21_ab_8__9_), .B(
        my_filter_first_coeff_mult_21_CARRYB_7__9_), .CI(
        my_filter_first_coeff_mult_21_SUMB_7__10_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_8__9_), .S(
        my_filter_first_coeff_mult_21_SUMB_8__9_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_8_8 ( .A(
        my_filter_first_coeff_mult_21_ab_8__8_), .B(
        my_filter_first_coeff_mult_21_CARRYB_7__8_), .CI(
        my_filter_first_coeff_mult_21_SUMB_7__9_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_8__8_), .S(
        my_filter_first_coeff_mult_21_SUMB_8__8_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_8_7 ( .A(
        my_filter_first_coeff_mult_21_ab_8__7_), .B(
        my_filter_first_coeff_mult_21_CARRYB_7__7_), .CI(
        my_filter_first_coeff_mult_21_SUMB_7__8_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_8__7_), .S(
        my_filter_first_coeff_mult_21_SUMB_8__7_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_8_6 ( .A(
        my_filter_first_coeff_mult_21_ab_8__6_), .B(
        my_filter_first_coeff_mult_21_CARRYB_7__6_), .CI(
        my_filter_first_coeff_mult_21_SUMB_7__7_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_8__6_), .S(
        my_filter_first_coeff_mult_21_SUMB_8__6_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_8_5 ( .A(
        my_filter_first_coeff_mult_21_ab_8__5_), .B(
        my_filter_first_coeff_mult_21_CARRYB_7__5_), .CI(
        my_filter_first_coeff_mult_21_SUMB_7__6_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_8__5_), .S(
        my_filter_first_coeff_mult_21_SUMB_8__5_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_8_4 ( .A(
        my_filter_first_coeff_mult_21_ab_8__4_), .B(
        my_filter_first_coeff_mult_21_CARRYB_7__4_), .CI(
        my_filter_first_coeff_mult_21_SUMB_7__5_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_8__4_), .S(
        my_filter_first_coeff_mult_21_SUMB_8__4_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_8_3 ( .A(
        my_filter_first_coeff_mult_21_ab_8__3_), .B(
        my_filter_first_coeff_mult_21_CARRYB_7__3_), .CI(
        my_filter_first_coeff_mult_21_SUMB_7__4_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_8__3_), .S(
        my_filter_first_coeff_mult_21_SUMB_8__3_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_8_2 ( .A(
        my_filter_first_coeff_mult_21_ab_8__2_), .B(
        my_filter_first_coeff_mult_21_CARRYB_7__2_), .CI(
        my_filter_first_coeff_mult_21_SUMB_7__3_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_8__2_), .S(
        my_filter_first_coeff_mult_21_SUMB_8__2_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_8_1 ( .A(
        my_filter_first_coeff_mult_21_ab_8__1_), .B(
        my_filter_first_coeff_mult_21_CARRYB_7__1_), .CI(
        my_filter_first_coeff_mult_21_SUMB_7__2_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_8__1_), .S(
        my_filter_first_coeff_mult_21_SUMB_8__1_) );
  FA_X1 my_filter_first_coeff_mult_21_S1_8_0 ( .A(
        my_filter_first_coeff_mult_21_ab_8__0_), .B(
        my_filter_first_coeff_mult_21_CARRYB_7__0_), .CI(
        my_filter_first_coeff_mult_21_SUMB_7__1_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_8__0_), .S(
        my_filter_first_coeff_mult_21_A1_6_) );
  FA_X1 my_filter_first_coeff_mult_21_S3_9_12 ( .A(
        my_filter_first_coeff_mult_21_ab_9__12_), .B(
        my_filter_first_coeff_mult_21_CARRYB_8__12_), .CI(
        my_filter_first_coeff_mult_21_ab_8__13_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_9__12_), .S(
        my_filter_first_coeff_mult_21_SUMB_9__12_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_9_11 ( .A(
        my_filter_first_coeff_mult_21_ab_9__11_), .B(
        my_filter_first_coeff_mult_21_CARRYB_8__11_), .CI(
        my_filter_first_coeff_mult_21_SUMB_8__12_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_9__11_), .S(
        my_filter_first_coeff_mult_21_SUMB_9__11_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_9_10 ( .A(
        my_filter_first_coeff_mult_21_ab_9__10_), .B(
        my_filter_first_coeff_mult_21_CARRYB_8__10_), .CI(
        my_filter_first_coeff_mult_21_SUMB_8__11_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_9__10_), .S(
        my_filter_first_coeff_mult_21_SUMB_9__10_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_9_9 ( .A(
        my_filter_first_coeff_mult_21_ab_9__9_), .B(
        my_filter_first_coeff_mult_21_CARRYB_8__9_), .CI(
        my_filter_first_coeff_mult_21_SUMB_8__10_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_9__9_), .S(
        my_filter_first_coeff_mult_21_SUMB_9__9_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_9_8 ( .A(
        my_filter_first_coeff_mult_21_ab_9__8_), .B(
        my_filter_first_coeff_mult_21_CARRYB_8__8_), .CI(
        my_filter_first_coeff_mult_21_SUMB_8__9_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_9__8_), .S(
        my_filter_first_coeff_mult_21_SUMB_9__8_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_9_7 ( .A(
        my_filter_first_coeff_mult_21_ab_9__7_), .B(
        my_filter_first_coeff_mult_21_CARRYB_8__7_), .CI(
        my_filter_first_coeff_mult_21_SUMB_8__8_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_9__7_), .S(
        my_filter_first_coeff_mult_21_SUMB_9__7_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_9_6 ( .A(
        my_filter_first_coeff_mult_21_ab_9__6_), .B(
        my_filter_first_coeff_mult_21_CARRYB_8__6_), .CI(
        my_filter_first_coeff_mult_21_SUMB_8__7_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_9__6_), .S(
        my_filter_first_coeff_mult_21_SUMB_9__6_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_9_5 ( .A(
        my_filter_first_coeff_mult_21_ab_9__5_), .B(
        my_filter_first_coeff_mult_21_CARRYB_8__5_), .CI(
        my_filter_first_coeff_mult_21_SUMB_8__6_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_9__5_), .S(
        my_filter_first_coeff_mult_21_SUMB_9__5_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_9_4 ( .A(
        my_filter_first_coeff_mult_21_ab_9__4_), .B(
        my_filter_first_coeff_mult_21_CARRYB_8__4_), .CI(
        my_filter_first_coeff_mult_21_SUMB_8__5_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_9__4_), .S(
        my_filter_first_coeff_mult_21_SUMB_9__4_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_9_3 ( .A(
        my_filter_first_coeff_mult_21_ab_9__3_), .B(
        my_filter_first_coeff_mult_21_CARRYB_8__3_), .CI(
        my_filter_first_coeff_mult_21_SUMB_8__4_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_9__3_), .S(
        my_filter_first_coeff_mult_21_SUMB_9__3_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_9_2 ( .A(
        my_filter_first_coeff_mult_21_ab_9__2_), .B(
        my_filter_first_coeff_mult_21_CARRYB_8__2_), .CI(
        my_filter_first_coeff_mult_21_SUMB_8__3_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_9__2_), .S(
        my_filter_first_coeff_mult_21_SUMB_9__2_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_9_1 ( .A(
        my_filter_first_coeff_mult_21_ab_9__1_), .B(
        my_filter_first_coeff_mult_21_CARRYB_8__1_), .CI(
        my_filter_first_coeff_mult_21_SUMB_8__2_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_9__1_), .S(
        my_filter_first_coeff_mult_21_SUMB_9__1_) );
  FA_X1 my_filter_first_coeff_mult_21_S1_9_0 ( .A(
        my_filter_first_coeff_mult_21_ab_9__0_), .B(
        my_filter_first_coeff_mult_21_CARRYB_8__0_), .CI(
        my_filter_first_coeff_mult_21_SUMB_8__1_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_9__0_), .S(
        my_filter_first_coeff_mult_21_A1_7_) );
  FA_X1 my_filter_first_coeff_mult_21_S3_10_12 ( .A(
        my_filter_first_coeff_mult_21_ab_10__12_), .B(
        my_filter_first_coeff_mult_21_CARRYB_9__12_), .CI(
        my_filter_first_coeff_mult_21_ab_9__13_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_10__12_), .S(
        my_filter_first_coeff_mult_21_SUMB_10__12_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_10_11 ( .A(
        my_filter_first_coeff_mult_21_ab_10__11_), .B(
        my_filter_first_coeff_mult_21_CARRYB_9__11_), .CI(
        my_filter_first_coeff_mult_21_SUMB_9__12_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_10__11_), .S(
        my_filter_first_coeff_mult_21_SUMB_10__11_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_10_10 ( .A(
        my_filter_first_coeff_mult_21_ab_10__10_), .B(
        my_filter_first_coeff_mult_21_CARRYB_9__10_), .CI(
        my_filter_first_coeff_mult_21_SUMB_9__11_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_10__10_), .S(
        my_filter_first_coeff_mult_21_SUMB_10__10_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_10_9 ( .A(
        my_filter_first_coeff_mult_21_ab_10__9_), .B(
        my_filter_first_coeff_mult_21_CARRYB_9__9_), .CI(
        my_filter_first_coeff_mult_21_SUMB_9__10_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_10__9_), .S(
        my_filter_first_coeff_mult_21_SUMB_10__9_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_10_8 ( .A(
        my_filter_first_coeff_mult_21_ab_10__8_), .B(
        my_filter_first_coeff_mult_21_CARRYB_9__8_), .CI(
        my_filter_first_coeff_mult_21_SUMB_9__9_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_10__8_), .S(
        my_filter_first_coeff_mult_21_SUMB_10__8_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_10_7 ( .A(
        my_filter_first_coeff_mult_21_ab_10__7_), .B(
        my_filter_first_coeff_mult_21_CARRYB_9__7_), .CI(
        my_filter_first_coeff_mult_21_SUMB_9__8_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_10__7_), .S(
        my_filter_first_coeff_mult_21_SUMB_10__7_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_10_6 ( .A(
        my_filter_first_coeff_mult_21_ab_10__6_), .B(
        my_filter_first_coeff_mult_21_CARRYB_9__6_), .CI(
        my_filter_first_coeff_mult_21_SUMB_9__7_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_10__6_), .S(
        my_filter_first_coeff_mult_21_SUMB_10__6_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_10_5 ( .A(
        my_filter_first_coeff_mult_21_ab_10__5_), .B(
        my_filter_first_coeff_mult_21_CARRYB_9__5_), .CI(
        my_filter_first_coeff_mult_21_SUMB_9__6_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_10__5_), .S(
        my_filter_first_coeff_mult_21_SUMB_10__5_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_10_4 ( .A(
        my_filter_first_coeff_mult_21_ab_10__4_), .B(
        my_filter_first_coeff_mult_21_CARRYB_9__4_), .CI(
        my_filter_first_coeff_mult_21_SUMB_9__5_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_10__4_), .S(
        my_filter_first_coeff_mult_21_SUMB_10__4_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_10_3 ( .A(
        my_filter_first_coeff_mult_21_ab_10__3_), .B(
        my_filter_first_coeff_mult_21_CARRYB_9__3_), .CI(
        my_filter_first_coeff_mult_21_SUMB_9__4_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_10__3_), .S(
        my_filter_first_coeff_mult_21_SUMB_10__3_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_10_2 ( .A(
        my_filter_first_coeff_mult_21_ab_10__2_), .B(
        my_filter_first_coeff_mult_21_CARRYB_9__2_), .CI(
        my_filter_first_coeff_mult_21_SUMB_9__3_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_10__2_), .S(
        my_filter_first_coeff_mult_21_SUMB_10__2_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_10_1 ( .A(
        my_filter_first_coeff_mult_21_ab_10__1_), .B(
        my_filter_first_coeff_mult_21_CARRYB_9__1_), .CI(
        my_filter_first_coeff_mult_21_SUMB_9__2_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_10__1_), .S(
        my_filter_first_coeff_mult_21_SUMB_10__1_) );
  FA_X1 my_filter_first_coeff_mult_21_S1_10_0 ( .A(
        my_filter_first_coeff_mult_21_ab_10__0_), .B(
        my_filter_first_coeff_mult_21_CARRYB_9__0_), .CI(
        my_filter_first_coeff_mult_21_SUMB_9__1_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_10__0_), .S(
        my_filter_first_coeff_mult_21_A1_8_) );
  FA_X1 my_filter_first_coeff_mult_21_S3_11_12 ( .A(
        my_filter_first_coeff_mult_21_ab_11__12_), .B(
        my_filter_first_coeff_mult_21_CARRYB_10__12_), .CI(
        my_filter_first_coeff_mult_21_ab_10__13_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_11__12_), .S(
        my_filter_first_coeff_mult_21_SUMB_11__12_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_11_11 ( .A(
        my_filter_first_coeff_mult_21_ab_11__11_), .B(
        my_filter_first_coeff_mult_21_CARRYB_10__11_), .CI(
        my_filter_first_coeff_mult_21_SUMB_10__12_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_11__11_), .S(
        my_filter_first_coeff_mult_21_SUMB_11__11_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_11_10 ( .A(
        my_filter_first_coeff_mult_21_ab_11__10_), .B(
        my_filter_first_coeff_mult_21_CARRYB_10__10_), .CI(
        my_filter_first_coeff_mult_21_SUMB_10__11_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_11__10_), .S(
        my_filter_first_coeff_mult_21_SUMB_11__10_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_11_9 ( .A(
        my_filter_first_coeff_mult_21_ab_11__9_), .B(
        my_filter_first_coeff_mult_21_CARRYB_10__9_), .CI(
        my_filter_first_coeff_mult_21_SUMB_10__10_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_11__9_), .S(
        my_filter_first_coeff_mult_21_SUMB_11__9_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_11_8 ( .A(
        my_filter_first_coeff_mult_21_ab_11__8_), .B(
        my_filter_first_coeff_mult_21_CARRYB_10__8_), .CI(
        my_filter_first_coeff_mult_21_SUMB_10__9_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_11__8_), .S(
        my_filter_first_coeff_mult_21_SUMB_11__8_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_11_7 ( .A(
        my_filter_first_coeff_mult_21_ab_11__7_), .B(
        my_filter_first_coeff_mult_21_CARRYB_10__7_), .CI(
        my_filter_first_coeff_mult_21_SUMB_10__8_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_11__7_), .S(
        my_filter_first_coeff_mult_21_SUMB_11__7_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_11_6 ( .A(
        my_filter_first_coeff_mult_21_ab_11__6_), .B(
        my_filter_first_coeff_mult_21_CARRYB_10__6_), .CI(
        my_filter_first_coeff_mult_21_SUMB_10__7_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_11__6_), .S(
        my_filter_first_coeff_mult_21_SUMB_11__6_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_11_5 ( .A(
        my_filter_first_coeff_mult_21_ab_11__5_), .B(
        my_filter_first_coeff_mult_21_CARRYB_10__5_), .CI(
        my_filter_first_coeff_mult_21_SUMB_10__6_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_11__5_), .S(
        my_filter_first_coeff_mult_21_SUMB_11__5_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_11_4 ( .A(
        my_filter_first_coeff_mult_21_ab_11__4_), .B(
        my_filter_first_coeff_mult_21_CARRYB_10__4_), .CI(
        my_filter_first_coeff_mult_21_SUMB_10__5_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_11__4_), .S(
        my_filter_first_coeff_mult_21_SUMB_11__4_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_11_3 ( .A(
        my_filter_first_coeff_mult_21_ab_11__3_), .B(
        my_filter_first_coeff_mult_21_CARRYB_10__3_), .CI(
        my_filter_first_coeff_mult_21_SUMB_10__4_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_11__3_), .S(
        my_filter_first_coeff_mult_21_SUMB_11__3_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_11_2 ( .A(
        my_filter_first_coeff_mult_21_ab_11__2_), .B(
        my_filter_first_coeff_mult_21_CARRYB_10__2_), .CI(
        my_filter_first_coeff_mult_21_SUMB_10__3_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_11__2_), .S(
        my_filter_first_coeff_mult_21_SUMB_11__2_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_11_1 ( .A(
        my_filter_first_coeff_mult_21_ab_11__1_), .B(
        my_filter_first_coeff_mult_21_CARRYB_10__1_), .CI(
        my_filter_first_coeff_mult_21_SUMB_10__2_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_11__1_), .S(
        my_filter_first_coeff_mult_21_SUMB_11__1_) );
  FA_X1 my_filter_first_coeff_mult_21_S1_11_0 ( .A(
        my_filter_first_coeff_mult_21_ab_11__0_), .B(
        my_filter_first_coeff_mult_21_CARRYB_10__0_), .CI(
        my_filter_first_coeff_mult_21_SUMB_10__1_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_11__0_), .S(
        my_filter_first_coeff_mult_21_A1_9_) );
  FA_X1 my_filter_first_coeff_mult_21_S3_12_12 ( .A(
        my_filter_first_coeff_mult_21_ab_12__12_), .B(
        my_filter_first_coeff_mult_21_CARRYB_11__12_), .CI(
        my_filter_first_coeff_mult_21_ab_11__13_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_12__12_), .S(
        my_filter_first_coeff_mult_21_SUMB_12__12_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_12_11 ( .A(
        my_filter_first_coeff_mult_21_ab_12__11_), .B(
        my_filter_first_coeff_mult_21_CARRYB_11__11_), .CI(
        my_filter_first_coeff_mult_21_SUMB_11__12_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_12__11_), .S(
        my_filter_first_coeff_mult_21_SUMB_12__11_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_12_10 ( .A(
        my_filter_first_coeff_mult_21_ab_12__10_), .B(
        my_filter_first_coeff_mult_21_CARRYB_11__10_), .CI(
        my_filter_first_coeff_mult_21_SUMB_11__11_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_12__10_), .S(
        my_filter_first_coeff_mult_21_SUMB_12__10_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_12_9 ( .A(
        my_filter_first_coeff_mult_21_ab_12__9_), .B(
        my_filter_first_coeff_mult_21_CARRYB_11__9_), .CI(
        my_filter_first_coeff_mult_21_SUMB_11__10_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_12__9_), .S(
        my_filter_first_coeff_mult_21_SUMB_12__9_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_12_8 ( .A(
        my_filter_first_coeff_mult_21_ab_12__8_), .B(
        my_filter_first_coeff_mult_21_CARRYB_11__8_), .CI(
        my_filter_first_coeff_mult_21_SUMB_11__9_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_12__8_), .S(
        my_filter_first_coeff_mult_21_SUMB_12__8_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_12_7 ( .A(
        my_filter_first_coeff_mult_21_ab_12__7_), .B(
        my_filter_first_coeff_mult_21_CARRYB_11__7_), .CI(
        my_filter_first_coeff_mult_21_SUMB_11__8_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_12__7_), .S(
        my_filter_first_coeff_mult_21_SUMB_12__7_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_12_6 ( .A(
        my_filter_first_coeff_mult_21_ab_12__6_), .B(
        my_filter_first_coeff_mult_21_CARRYB_11__6_), .CI(
        my_filter_first_coeff_mult_21_SUMB_11__7_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_12__6_), .S(
        my_filter_first_coeff_mult_21_SUMB_12__6_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_12_5 ( .A(
        my_filter_first_coeff_mult_21_ab_12__5_), .B(
        my_filter_first_coeff_mult_21_CARRYB_11__5_), .CI(
        my_filter_first_coeff_mult_21_SUMB_11__6_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_12__5_), .S(
        my_filter_first_coeff_mult_21_SUMB_12__5_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_12_4 ( .A(
        my_filter_first_coeff_mult_21_ab_12__4_), .B(
        my_filter_first_coeff_mult_21_CARRYB_11__4_), .CI(
        my_filter_first_coeff_mult_21_SUMB_11__5_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_12__4_), .S(
        my_filter_first_coeff_mult_21_SUMB_12__4_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_12_3 ( .A(
        my_filter_first_coeff_mult_21_ab_12__3_), .B(
        my_filter_first_coeff_mult_21_CARRYB_11__3_), .CI(
        my_filter_first_coeff_mult_21_SUMB_11__4_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_12__3_), .S(
        my_filter_first_coeff_mult_21_SUMB_12__3_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_12_2 ( .A(
        my_filter_first_coeff_mult_21_ab_12__2_), .B(
        my_filter_first_coeff_mult_21_CARRYB_11__2_), .CI(
        my_filter_first_coeff_mult_21_SUMB_11__3_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_12__2_), .S(
        my_filter_first_coeff_mult_21_SUMB_12__2_) );
  FA_X1 my_filter_first_coeff_mult_21_S2_12_1 ( .A(
        my_filter_first_coeff_mult_21_ab_12__1_), .B(
        my_filter_first_coeff_mult_21_CARRYB_11__1_), .CI(
        my_filter_first_coeff_mult_21_SUMB_11__2_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_12__1_), .S(
        my_filter_first_coeff_mult_21_SUMB_12__1_) );
  FA_X1 my_filter_first_coeff_mult_21_S1_12_0 ( .A(
        my_filter_first_coeff_mult_21_ab_12__0_), .B(
        my_filter_first_coeff_mult_21_CARRYB_11__0_), .CI(
        my_filter_first_coeff_mult_21_SUMB_11__1_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_12__0_), .S(
        my_filter_first_coeff_mult_21_A1_10_) );
  FA_X1 my_filter_first_coeff_mult_21_S14_13 ( .A(
        my_filter_first_coeff_mult_21_n100), .B(
        my_filter_first_coeff_mult_21_n86), .CI(
        my_filter_first_coeff_mult_21_ab_13__13_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_13__13_), .S(
        my_filter_first_coeff_mult_21_SUMB_13__13_) );
  FA_X1 my_filter_first_coeff_mult_21_S5_12 ( .A(
        my_filter_first_coeff_mult_21_ab_13__12_), .B(
        my_filter_first_coeff_mult_21_CARRYB_12__12_), .CI(
        my_filter_first_coeff_mult_21_ab_12__13_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_13__12_), .S(
        my_filter_first_coeff_mult_21_SUMB_13__12_) );
  FA_X1 my_filter_first_coeff_mult_21_S4_11 ( .A(
        my_filter_first_coeff_mult_21_ab_13__11_), .B(
        my_filter_first_coeff_mult_21_CARRYB_12__11_), .CI(
        my_filter_first_coeff_mult_21_SUMB_12__12_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_13__11_), .S(
        my_filter_first_coeff_mult_21_SUMB_13__11_) );
  FA_X1 my_filter_first_coeff_mult_21_S4_10 ( .A(
        my_filter_first_coeff_mult_21_ab_13__10_), .B(
        my_filter_first_coeff_mult_21_CARRYB_12__10_), .CI(
        my_filter_first_coeff_mult_21_SUMB_12__11_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_13__10_), .S(
        my_filter_first_coeff_mult_21_SUMB_13__10_) );
  FA_X1 my_filter_first_coeff_mult_21_S4_9 ( .A(
        my_filter_first_coeff_mult_21_ab_13__9_), .B(
        my_filter_first_coeff_mult_21_CARRYB_12__9_), .CI(
        my_filter_first_coeff_mult_21_SUMB_12__10_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_13__9_), .S(
        my_filter_first_coeff_mult_21_SUMB_13__9_) );
  FA_X1 my_filter_first_coeff_mult_21_S4_8 ( .A(
        my_filter_first_coeff_mult_21_ab_13__8_), .B(
        my_filter_first_coeff_mult_21_CARRYB_12__8_), .CI(
        my_filter_first_coeff_mult_21_SUMB_12__9_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_13__8_), .S(
        my_filter_first_coeff_mult_21_SUMB_13__8_) );
  FA_X1 my_filter_first_coeff_mult_21_S4_7 ( .A(
        my_filter_first_coeff_mult_21_ab_13__7_), .B(
        my_filter_first_coeff_mult_21_CARRYB_12__7_), .CI(
        my_filter_first_coeff_mult_21_SUMB_12__8_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_13__7_), .S(
        my_filter_first_coeff_mult_21_SUMB_13__7_) );
  FA_X1 my_filter_first_coeff_mult_21_S4_6 ( .A(
        my_filter_first_coeff_mult_21_ab_13__6_), .B(
        my_filter_first_coeff_mult_21_CARRYB_12__6_), .CI(
        my_filter_first_coeff_mult_21_SUMB_12__7_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_13__6_), .S(
        my_filter_first_coeff_mult_21_SUMB_13__6_) );
  FA_X1 my_filter_first_coeff_mult_21_S4_5 ( .A(
        my_filter_first_coeff_mult_21_ab_13__5_), .B(
        my_filter_first_coeff_mult_21_CARRYB_12__5_), .CI(
        my_filter_first_coeff_mult_21_SUMB_12__6_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_13__5_), .S(
        my_filter_first_coeff_mult_21_SUMB_13__5_) );
  FA_X1 my_filter_first_coeff_mult_21_S4_4 ( .A(
        my_filter_first_coeff_mult_21_ab_13__4_), .B(
        my_filter_first_coeff_mult_21_CARRYB_12__4_), .CI(
        my_filter_first_coeff_mult_21_SUMB_12__5_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_13__4_), .S(
        my_filter_first_coeff_mult_21_SUMB_13__4_) );
  FA_X1 my_filter_first_coeff_mult_21_S4_3 ( .A(
        my_filter_first_coeff_mult_21_ab_13__3_), .B(
        my_filter_first_coeff_mult_21_CARRYB_12__3_), .CI(
        my_filter_first_coeff_mult_21_SUMB_12__4_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_13__3_), .S(
        my_filter_first_coeff_mult_21_SUMB_13__3_) );
  FA_X1 my_filter_first_coeff_mult_21_S4_2 ( .A(
        my_filter_first_coeff_mult_21_ab_13__2_), .B(
        my_filter_first_coeff_mult_21_CARRYB_12__2_), .CI(
        my_filter_first_coeff_mult_21_SUMB_12__3_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_13__2_), .S(
        my_filter_first_coeff_mult_21_SUMB_13__2_) );
  FA_X1 my_filter_first_coeff_mult_21_S4_1 ( .A(
        my_filter_first_coeff_mult_21_ab_13__1_), .B(
        my_filter_first_coeff_mult_21_CARRYB_12__1_), .CI(
        my_filter_first_coeff_mult_21_SUMB_12__2_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_13__1_), .S(
        my_filter_first_coeff_mult_21_SUMB_13__1_) );
  FA_X1 my_filter_first_coeff_mult_21_S4_0 ( .A(
        my_filter_first_coeff_mult_21_ab_13__0_), .B(
        my_filter_first_coeff_mult_21_CARRYB_12__0_), .CI(
        my_filter_first_coeff_mult_21_SUMB_12__1_), .CO(
        my_filter_first_coeff_mult_21_CARRYB_13__0_), .S(
        my_filter_first_coeff_mult_21_SUMB_13__0_) );
  FA_X1 my_filter_first_coeff_mult_21_S14_13_0 ( .A(my_filter_q_reg_samp_13_), 
        .B(my_filter_q_reg_coeff[153]), .CI(
        my_filter_first_coeff_mult_21_SUMB_13__0_), .CO(
        my_filter_first_coeff_mult_21_A2_12_), .S(my_filter_data_sum[140]) );
  NAND2_X1 my_filter_first_coeff_mult_21_FS_1_U72 ( .A1(
        my_filter_first_coeff_mult_21_A2_12_), .A2(
        my_filter_first_coeff_mult_21_n29), .ZN(
        my_filter_first_coeff_mult_21_FS_1_n56) );
  INV_X1 my_filter_first_coeff_mult_21_FS_1_U71 ( .A(
        my_filter_first_coeff_mult_21_FS_1_n59), .ZN(my_filter_data_sum[141])
         );
  OAI21_X1 my_filter_first_coeff_mult_21_FS_1_U70 ( .B1(
        my_filter_first_coeff_mult_21_A2_12_), .B2(
        my_filter_first_coeff_mult_21_n29), .A(
        my_filter_first_coeff_mult_21_FS_1_n56), .ZN(
        my_filter_first_coeff_mult_21_FS_1_n59) );
  AND2_X1 my_filter_first_coeff_mult_21_FS_1_U69 ( .A1(
        my_filter_first_coeff_mult_21_n52), .A2(
        my_filter_first_coeff_mult_21_n50), .ZN(
        my_filter_first_coeff_mult_21_FS_1_n20) );
  AND2_X1 my_filter_first_coeff_mult_21_FS_1_U68 ( .A1(
        my_filter_first_coeff_mult_21_n51), .A2(
        my_filter_first_coeff_mult_21_n46), .ZN(
        my_filter_first_coeff_mult_21_FS_1_n28) );
  NAND2_X1 my_filter_first_coeff_mult_21_FS_1_U66 ( .A1(
        my_filter_first_coeff_mult_21_n48), .A2(
        my_filter_first_coeff_mult_21_n47), .ZN(
        my_filter_first_coeff_mult_21_FS_1_n17) );
  NAND2_X1 my_filter_first_coeff_mult_21_FS_1_U65 ( .A1(
        my_filter_first_coeff_mult_21_n49), .A2(
        my_filter_first_coeff_mult_21_n45), .ZN(
        my_filter_first_coeff_mult_21_FS_1_n25) );
  NOR2_X1 my_filter_first_coeff_mult_21_FS_1_U64 ( .A1(
        my_filter_first_coeff_mult_21_n48), .A2(
        my_filter_first_coeff_mult_21_n47), .ZN(
        my_filter_first_coeff_mult_21_FS_1_n15) );
  NOR2_X1 my_filter_first_coeff_mult_21_FS_1_U63 ( .A1(
        my_filter_first_coeff_mult_21_n49), .A2(
        my_filter_first_coeff_mult_21_n45), .ZN(
        my_filter_first_coeff_mult_21_FS_1_n23) );
  NOR2_X1 my_filter_first_coeff_mult_21_FS_1_U61 ( .A1(
        my_filter_first_coeff_mult_21_n52), .A2(
        my_filter_first_coeff_mult_21_n50), .ZN(
        my_filter_first_coeff_mult_21_FS_1_n21) );
  NOR2_X1 my_filter_first_coeff_mult_21_FS_1_U60 ( .A1(
        my_filter_first_coeff_mult_21_n51), .A2(
        my_filter_first_coeff_mult_21_n46), .ZN(
        my_filter_first_coeff_mult_21_FS_1_n29) );
  AND2_X1 my_filter_first_coeff_mult_21_FS_1_U59 ( .A1(
        my_filter_first_coeff_mult_21_n43), .A2(
        my_filter_first_coeff_mult_21_n33), .ZN(
        my_filter_first_coeff_mult_21_FS_1_n36) );
  AND2_X1 my_filter_first_coeff_mult_21_FS_1_U58 ( .A1(
        my_filter_first_coeff_mult_21_n34), .A2(
        my_filter_first_coeff_mult_21_n31), .ZN(
        my_filter_first_coeff_mult_21_FS_1_n44) );
  AND2_X1 my_filter_first_coeff_mult_21_FS_1_U56 ( .A1(
        my_filter_first_coeff_mult_21_n42), .A2(
        my_filter_first_coeff_mult_21_n30), .ZN(
        my_filter_first_coeff_mult_21_FS_1_n52) );
  NAND2_X1 my_filter_first_coeff_mult_21_FS_1_U55 ( .A1(
        my_filter_first_coeff_mult_21_n41), .A2(
        my_filter_first_coeff_mult_21_n32), .ZN(
        my_filter_first_coeff_mult_21_FS_1_n33) );
  NAND2_X1 my_filter_first_coeff_mult_21_FS_1_U54 ( .A1(
        my_filter_first_coeff_mult_21_n40), .A2(
        my_filter_first_coeff_mult_21_n37), .ZN(
        my_filter_first_coeff_mult_21_FS_1_n41) );
  NAND2_X1 my_filter_first_coeff_mult_21_FS_1_U53 ( .A1(
        my_filter_first_coeff_mult_21_n39), .A2(
        my_filter_first_coeff_mult_21_n36), .ZN(
        my_filter_first_coeff_mult_21_FS_1_n49) );
  NAND2_X1 my_filter_first_coeff_mult_21_FS_1_U51 ( .A1(
        my_filter_first_coeff_mult_21_n38), .A2(
        my_filter_first_coeff_mult_21_n35), .ZN(
        my_filter_first_coeff_mult_21_FS_1_n57) );
  NAND2_X1 my_filter_first_coeff_mult_21_FS_1_U50 ( .A1(
        my_filter_first_coeff_mult_21_FS_1_n70), .A2(
        my_filter_first_coeff_mult_21_FS_1_n57), .ZN(
        my_filter_first_coeff_mult_21_FS_1_n58) );
  NOR2_X1 my_filter_first_coeff_mult_21_FS_1_U49 ( .A1(
        my_filter_first_coeff_mult_21_n41), .A2(
        my_filter_first_coeff_mult_21_n32), .ZN(
        my_filter_first_coeff_mult_21_FS_1_n31) );
  NOR2_X1 my_filter_first_coeff_mult_21_FS_1_U48 ( .A1(
        my_filter_first_coeff_mult_21_n40), .A2(
        my_filter_first_coeff_mult_21_n37), .ZN(
        my_filter_first_coeff_mult_21_FS_1_n39) );
  NOR2_X1 my_filter_first_coeff_mult_21_FS_1_U46 ( .A1(
        my_filter_first_coeff_mult_21_n39), .A2(
        my_filter_first_coeff_mult_21_n36), .ZN(
        my_filter_first_coeff_mult_21_FS_1_n47) );
  NOR2_X1 my_filter_first_coeff_mult_21_FS_1_U45 ( .A1(
        my_filter_first_coeff_mult_21_n38), .A2(
        my_filter_first_coeff_mult_21_n35), .ZN(
        my_filter_first_coeff_mult_21_FS_1_n55) );
  NOR2_X1 my_filter_first_coeff_mult_21_FS_1_U44 ( .A1(
        my_filter_first_coeff_mult_21_n43), .A2(
        my_filter_first_coeff_mult_21_n33), .ZN(
        my_filter_first_coeff_mult_21_FS_1_n37) );
  NOR2_X1 my_filter_first_coeff_mult_21_FS_1_U43 ( .A1(
        my_filter_first_coeff_mult_21_n34), .A2(
        my_filter_first_coeff_mult_21_n31), .ZN(
        my_filter_first_coeff_mult_21_FS_1_n45) );
  NOR2_X1 my_filter_first_coeff_mult_21_FS_1_U41 ( .A1(
        my_filter_first_coeff_mult_21_n42), .A2(
        my_filter_first_coeff_mult_21_n30), .ZN(
        my_filter_first_coeff_mult_21_FS_1_n53) );
  OAI21_X1 my_filter_first_coeff_mult_21_FS_1_U40 ( .B1(
        my_filter_first_coeff_mult_21_FS_1_n55), .B2(
        my_filter_first_coeff_mult_21_FS_1_n56), .A(
        my_filter_first_coeff_mult_21_FS_1_n57), .ZN(
        my_filter_first_coeff_mult_21_FS_1_n51) );
  INV_X1 my_filter_first_coeff_mult_21_FS_1_U39 ( .A(
        my_filter_first_coeff_mult_21_FS_1_n15), .ZN(
        my_filter_first_coeff_mult_21_FS_1_n60) );
  NAND2_X1 my_filter_first_coeff_mult_21_FS_1_U38 ( .A1(
        my_filter_first_coeff_mult_21_FS_1_n60), .A2(
        my_filter_first_coeff_mult_21_FS_1_n17), .ZN(
        my_filter_first_coeff_mult_21_FS_1_n18) );
  INV_X1 my_filter_first_coeff_mult_21_FS_1_U36 ( .A(
        my_filter_first_coeff_mult_21_FS_1_n23), .ZN(
        my_filter_first_coeff_mult_21_FS_1_n62) );
  NAND2_X1 my_filter_first_coeff_mult_21_FS_1_U35 ( .A1(
        my_filter_first_coeff_mult_21_FS_1_n62), .A2(
        my_filter_first_coeff_mult_21_FS_1_n25), .ZN(
        my_filter_first_coeff_mult_21_FS_1_n26) );
  NOR2_X1 my_filter_first_coeff_mult_21_FS_1_U34 ( .A1(
        my_filter_first_coeff_mult_21_FS_1_n20), .A2(
        my_filter_first_coeff_mult_21_FS_1_n21), .ZN(
        my_filter_first_coeff_mult_21_FS_1_n22) );
  NOR2_X1 my_filter_first_coeff_mult_21_FS_1_U33 ( .A1(
        my_filter_first_coeff_mult_21_FS_1_n28), .A2(
        my_filter_first_coeff_mult_21_FS_1_n29), .ZN(
        my_filter_first_coeff_mult_21_FS_1_n30) );
  INV_X1 my_filter_first_coeff_mult_21_FS_1_U31 ( .A(
        my_filter_first_coeff_mult_21_FS_1_n39), .ZN(
        my_filter_first_coeff_mult_21_FS_1_n66) );
  INV_X1 my_filter_first_coeff_mult_21_FS_1_U30 ( .A(
        my_filter_first_coeff_mult_21_FS_1_n47), .ZN(
        my_filter_first_coeff_mult_21_FS_1_n68) );
  INV_X1 my_filter_first_coeff_mult_21_FS_1_U29 ( .A(
        my_filter_first_coeff_mult_21_FS_1_n55), .ZN(
        my_filter_first_coeff_mult_21_FS_1_n70) );
  INV_X1 my_filter_first_coeff_mult_21_FS_1_U28 ( .A(
        my_filter_first_coeff_mult_21_FS_1_n31), .ZN(
        my_filter_first_coeff_mult_21_FS_1_n64) );
  NAND2_X1 my_filter_first_coeff_mult_21_FS_1_U26 ( .A1(
        my_filter_first_coeff_mult_21_FS_1_n64), .A2(
        my_filter_first_coeff_mult_21_FS_1_n33), .ZN(
        my_filter_first_coeff_mult_21_FS_1_n34) );
  NOR2_X1 my_filter_first_coeff_mult_21_FS_1_U25 ( .A1(
        my_filter_first_coeff_mult_21_FS_1_n36), .A2(
        my_filter_first_coeff_mult_21_FS_1_n37), .ZN(
        my_filter_first_coeff_mult_21_FS_1_n38) );
  NOR2_X1 my_filter_first_coeff_mult_21_FS_1_U24 ( .A1(
        my_filter_first_coeff_mult_21_FS_1_n44), .A2(
        my_filter_first_coeff_mult_21_FS_1_n45), .ZN(
        my_filter_first_coeff_mult_21_FS_1_n46) );
  NOR2_X1 my_filter_first_coeff_mult_21_FS_1_U23 ( .A1(
        my_filter_first_coeff_mult_21_FS_1_n52), .A2(
        my_filter_first_coeff_mult_21_FS_1_n53), .ZN(
        my_filter_first_coeff_mult_21_FS_1_n54) );
  NAND2_X1 my_filter_first_coeff_mult_21_FS_1_U21 ( .A1(
        my_filter_first_coeff_mult_21_FS_1_n66), .A2(
        my_filter_first_coeff_mult_21_FS_1_n41), .ZN(
        my_filter_first_coeff_mult_21_FS_1_n42) );
  NAND2_X1 my_filter_first_coeff_mult_21_FS_1_U20 ( .A1(
        my_filter_first_coeff_mult_21_FS_1_n68), .A2(
        my_filter_first_coeff_mult_21_FS_1_n49), .ZN(
        my_filter_first_coeff_mult_21_FS_1_n50) );
  OAI21_X1 my_filter_first_coeff_mult_21_FS_1_U19 ( .B1(
        my_filter_first_coeff_mult_21_FS_1_n15), .B2(
        my_filter_first_coeff_mult_21_FS_1_n16), .A(
        my_filter_first_coeff_mult_21_FS_1_n17), .ZN(
        my_filter_first_coeff_mult_21_FS_1_n13) );
  OAI21_X1 my_filter_first_coeff_mult_21_FS_1_U18 ( .B1(
        my_filter_first_coeff_mult_21_FS_1_n23), .B2(
        my_filter_first_coeff_mult_21_FS_1_n24), .A(
        my_filter_first_coeff_mult_21_FS_1_n25), .ZN(
        my_filter_first_coeff_mult_21_FS_1_n19) );
  OAI21_X1 my_filter_first_coeff_mult_21_FS_1_U16 ( .B1(
        my_filter_first_coeff_mult_21_FS_1_n31), .B2(
        my_filter_first_coeff_mult_21_FS_1_n32), .A(
        my_filter_first_coeff_mult_21_FS_1_n33), .ZN(
        my_filter_first_coeff_mult_21_FS_1_n27) );
  OAI21_X1 my_filter_first_coeff_mult_21_FS_1_U13 ( .B1(
        my_filter_first_coeff_mult_21_FS_1_n39), .B2(
        my_filter_first_coeff_mult_21_FS_1_n40), .A(
        my_filter_first_coeff_mult_21_FS_1_n41), .ZN(
        my_filter_first_coeff_mult_21_FS_1_n35) );
  OAI21_X1 my_filter_first_coeff_mult_21_FS_1_U12 ( .B1(
        my_filter_first_coeff_mult_21_FS_1_n47), .B2(
        my_filter_first_coeff_mult_21_FS_1_n48), .A(
        my_filter_first_coeff_mult_21_FS_1_n49), .ZN(
        my_filter_first_coeff_mult_21_FS_1_n43) );
  INV_X1 my_filter_first_coeff_mult_21_FS_1_U11 ( .A(
        my_filter_first_coeff_mult_21_FS_1_n21), .ZN(
        my_filter_first_coeff_mult_21_FS_1_n61) );
  AOI21_X1 my_filter_first_coeff_mult_21_FS_1_U10 ( .B1(
        my_filter_first_coeff_mult_21_FS_1_n61), .B2(
        my_filter_first_coeff_mult_21_FS_1_n19), .A(
        my_filter_first_coeff_mult_21_FS_1_n20), .ZN(
        my_filter_first_coeff_mult_21_FS_1_n16) );
  INV_X1 my_filter_first_coeff_mult_21_FS_1_U9 ( .A(
        my_filter_first_coeff_mult_21_FS_1_n29), .ZN(
        my_filter_first_coeff_mult_21_FS_1_n63) );
  AOI21_X1 my_filter_first_coeff_mult_21_FS_1_U8 ( .B1(
        my_filter_first_coeff_mult_21_FS_1_n63), .B2(
        my_filter_first_coeff_mult_21_FS_1_n27), .A(
        my_filter_first_coeff_mult_21_FS_1_n28), .ZN(
        my_filter_first_coeff_mult_21_FS_1_n24) );
  INV_X1 my_filter_first_coeff_mult_21_FS_1_U7 ( .A(
        my_filter_first_coeff_mult_21_FS_1_n37), .ZN(
        my_filter_first_coeff_mult_21_FS_1_n65) );
  AOI21_X1 my_filter_first_coeff_mult_21_FS_1_U6 ( .B1(
        my_filter_first_coeff_mult_21_FS_1_n65), .B2(
        my_filter_first_coeff_mult_21_FS_1_n35), .A(
        my_filter_first_coeff_mult_21_FS_1_n36), .ZN(
        my_filter_first_coeff_mult_21_FS_1_n32) );
  INV_X1 my_filter_first_coeff_mult_21_FS_1_U5 ( .A(
        my_filter_first_coeff_mult_21_FS_1_n45), .ZN(
        my_filter_first_coeff_mult_21_FS_1_n67) );
  AOI21_X1 my_filter_first_coeff_mult_21_FS_1_U4 ( .B1(
        my_filter_first_coeff_mult_21_FS_1_n67), .B2(
        my_filter_first_coeff_mult_21_FS_1_n43), .A(
        my_filter_first_coeff_mult_21_FS_1_n44), .ZN(
        my_filter_first_coeff_mult_21_FS_1_n40) );
  INV_X1 my_filter_first_coeff_mult_21_FS_1_U3 ( .A(
        my_filter_first_coeff_mult_21_FS_1_n53), .ZN(
        my_filter_first_coeff_mult_21_FS_1_n69) );
  AOI21_X1 my_filter_first_coeff_mult_21_FS_1_U2 ( .B1(
        my_filter_first_coeff_mult_21_FS_1_n69), .B2(
        my_filter_first_coeff_mult_21_FS_1_n51), .A(
        my_filter_first_coeff_mult_21_FS_1_n52), .ZN(
        my_filter_first_coeff_mult_21_FS_1_n48) );
  XOR2_X1 my_filter_first_coeff_mult_21_FS_1_U67 ( .A(
        my_filter_first_coeff_mult_21_FS_1_n56), .B(
        my_filter_first_coeff_mult_21_FS_1_n58), .Z(my_filter_data_sum[142])
         );
  XOR2_X1 my_filter_first_coeff_mult_21_FS_1_U62 ( .A(
        my_filter_first_coeff_mult_21_FS_1_n51), .B(
        my_filter_first_coeff_mult_21_FS_1_n54), .Z(my_filter_data_sum[143])
         );
  XOR2_X1 my_filter_first_coeff_mult_21_FS_1_U57 ( .A(
        my_filter_first_coeff_mult_21_FS_1_n50), .B(
        my_filter_first_coeff_mult_21_FS_1_n48), .Z(my_filter_data_sum[144])
         );
  XOR2_X1 my_filter_first_coeff_mult_21_FS_1_U52 ( .A(
        my_filter_first_coeff_mult_21_FS_1_n43), .B(
        my_filter_first_coeff_mult_21_FS_1_n46), .Z(my_filter_data_sum[145])
         );
  XOR2_X1 my_filter_first_coeff_mult_21_FS_1_U47 ( .A(
        my_filter_first_coeff_mult_21_FS_1_n42), .B(
        my_filter_first_coeff_mult_21_FS_1_n40), .Z(my_filter_data_sum[146])
         );
  XOR2_X1 my_filter_first_coeff_mult_21_FS_1_U42 ( .A(
        my_filter_first_coeff_mult_21_FS_1_n35), .B(
        my_filter_first_coeff_mult_21_FS_1_n38), .Z(my_filter_data_sum[147])
         );
  XOR2_X1 my_filter_first_coeff_mult_21_FS_1_U37 ( .A(
        my_filter_first_coeff_mult_21_FS_1_n34), .B(
        my_filter_first_coeff_mult_21_FS_1_n32), .Z(my_filter_data_sum[148])
         );
  XOR2_X1 my_filter_first_coeff_mult_21_FS_1_U32 ( .A(
        my_filter_first_coeff_mult_21_FS_1_n27), .B(
        my_filter_first_coeff_mult_21_FS_1_n30), .Z(my_filter_data_sum[149])
         );
  XOR2_X1 my_filter_first_coeff_mult_21_FS_1_U27 ( .A(
        my_filter_first_coeff_mult_21_FS_1_n26), .B(
        my_filter_first_coeff_mult_21_FS_1_n24), .Z(my_filter_data_sum[150])
         );
  XOR2_X1 my_filter_first_coeff_mult_21_FS_1_U22 ( .A(
        my_filter_first_coeff_mult_21_FS_1_n19), .B(
        my_filter_first_coeff_mult_21_FS_1_n22), .Z(my_filter_data_sum[151])
         );
  XOR2_X1 my_filter_first_coeff_mult_21_FS_1_U17 ( .A(
        my_filter_first_coeff_mult_21_FS_1_n18), .B(
        my_filter_first_coeff_mult_21_FS_1_n16), .Z(my_filter_data_sum[152])
         );
  XOR2_X1 my_filter_first_coeff_mult_21_FS_1_U15 ( .A(
        my_filter_first_coeff_mult_21_n27), .B(
        my_filter_first_coeff_mult_21_n44), .Z(
        my_filter_first_coeff_mult_21_FS_1_n14) );
  XOR2_X1 my_filter_first_coeff_mult_21_FS_1_U14 ( .A(
        my_filter_first_coeff_mult_21_FS_1_n13), .B(
        my_filter_first_coeff_mult_21_FS_1_n14), .Z(my_filter_data_sum[153])
         );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U276 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_12__12_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U275 ( .A1(
        my_filter_q_reg_chain_1__11_), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_11__13_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U274 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_11__12_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U273 ( .A1(
        my_filter_q_reg_chain_1__10_), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_10__13_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U272 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_10__12_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U271 ( .A1(
        my_filter_q_reg_chain_1__9_), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_9__13_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U270 ( .A1(
        my_filter_q_reg_coeff[136]), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_13__10_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U269 ( .A1(
        my_filter_q_reg_coeff[137]), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_13__11_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U268 ( .A1(
        my_filter_q_reg_coeff[135]), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_13__9_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U267 ( .A1(
        my_filter_q_reg_coeff[138]), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_13__12_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U266 ( .A1(
        my_filter_q_reg_chain_1__12_), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_12__13_) );
  INV_X1 my_filter_adder_mult_0_multiplication_mult_21_U265 ( .A(
        my_filter_q_reg_chain_1__9_), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_n90) );
  INV_X1 my_filter_adder_mult_0_multiplication_mult_21_U264 ( .A(
        my_filter_q_reg_chain_1__12_), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_n87) );
  INV_X1 my_filter_adder_mult_0_multiplication_mult_21_U263 ( .A(
        my_filter_q_reg_chain_1__11_), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_n88) );
  INV_X1 my_filter_adder_mult_0_multiplication_mult_21_U262 ( .A(
        my_filter_q_reg_chain_1__10_), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_n89) );
  INV_X1 my_filter_adder_mult_0_multiplication_mult_21_U261 ( .A(
        my_filter_q_reg_chain_1__8_), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_n91) );
  INV_X1 my_filter_adder_mult_0_multiplication_mult_21_U260 ( .A(
        my_filter_q_reg_chain_1__13_), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_n86) );
  AND2_X1 my_filter_adder_mult_0_multiplication_mult_21_U259 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_ab_0__13_), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_ab_1__12_), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_n15) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U258 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_2__12_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U257 ( .A1(
        my_filter_q_reg_chain_1__1_), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_1__13_) );
  AND3_X1 my_filter_adder_mult_0_multiplication_mult_21_U256 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_ab_1__1_), .A2(
        my_filter_q_reg_coeff[126]), .A3(my_filter_q_reg_chain_1__0_), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_1__0_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U255 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_12__0_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U254 ( .A1(
        my_filter_q_reg_coeff[126]), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_13__0_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U253 ( .A1(
        my_filter_q_reg_chain_1__8_), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_8__13_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U252 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n101), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_9__12_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U251 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_8__12_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U250 ( .A1(
        my_filter_q_reg_chain_1__7_), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_7__13_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U249 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_7__12_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U248 ( .A1(
        my_filter_q_reg_chain_1__6_), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_6__13_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U247 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_6__12_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U246 ( .A1(
        my_filter_q_reg_chain_1__5_), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_5__13_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U245 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_5__12_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U244 ( .A1(
        my_filter_q_reg_chain_1__4_), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_4__13_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U243 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_4__12_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U242 ( .A1(
        my_filter_q_reg_chain_1__3_), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_3__13_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U241 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_3__12_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U240 ( .A1(
        my_filter_q_reg_chain_1__2_), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_2__13_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U239 ( .A1(
        my_filter_q_reg_coeff[134]), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_13__8_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U238 ( .A1(
        my_filter_q_reg_coeff[132]), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_13__6_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U237 ( .A1(
        my_filter_q_reg_coeff[133]), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_13__7_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U236 ( .A1(
        my_filter_q_reg_coeff[130]), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_13__4_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U235 ( .A1(
        my_filter_q_reg_coeff[131]), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_13__5_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U234 ( .A1(
        my_filter_q_reg_coeff[128]), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_13__2_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U233 ( .A1(
        my_filter_q_reg_coeff[129]), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_13__3_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U232 ( .A1(
        my_filter_q_reg_coeff[127]), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_13__1_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U231 ( .A1(
        my_filter_q_reg_chain_1__0_), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_0__13_) );
  INV_X1 my_filter_adder_mult_0_multiplication_mult_21_U230 ( .A(
        my_filter_q_reg_coeff[139]), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_n100) );
  INV_X1 my_filter_adder_mult_0_multiplication_mult_21_U229 ( .A(
        my_filter_q_reg_coeff[126]), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_n113) );
  INV_X1 my_filter_adder_mult_0_multiplication_mult_21_U228 ( .A(
        my_filter_q_reg_chain_1__0_), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_n99) );
  INV_X1 my_filter_adder_mult_0_multiplication_mult_21_U227 ( .A(
        my_filter_q_reg_coeff[127]), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_n112) );
  INV_X1 my_filter_adder_mult_0_multiplication_mult_21_U226 ( .A(
        my_filter_q_reg_chain_1__1_), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_n98) );
  INV_X1 my_filter_adder_mult_0_multiplication_mult_21_U225 ( .A(
        my_filter_q_reg_coeff[138]), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_n101) );
  INV_X1 my_filter_adder_mult_0_multiplication_mult_21_U224 ( .A(
        my_filter_q_reg_coeff[136]), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_n103) );
  INV_X1 my_filter_adder_mult_0_multiplication_mult_21_U223 ( .A(
        my_filter_q_reg_coeff[137]), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_n102) );
  INV_X1 my_filter_adder_mult_0_multiplication_mult_21_U222 ( .A(
        my_filter_q_reg_coeff[134]), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_n105) );
  INV_X1 my_filter_adder_mult_0_multiplication_mult_21_U221 ( .A(
        my_filter_q_reg_coeff[135]), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_n104) );
  INV_X1 my_filter_adder_mult_0_multiplication_mult_21_U220 ( .A(
        my_filter_q_reg_coeff[132]), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_n107) );
  INV_X1 my_filter_adder_mult_0_multiplication_mult_21_U219 ( .A(
        my_filter_q_reg_coeff[133]), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_n106) );
  INV_X1 my_filter_adder_mult_0_multiplication_mult_21_U218 ( .A(
        my_filter_q_reg_coeff[128]), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_n111) );
  INV_X1 my_filter_adder_mult_0_multiplication_mult_21_U217 ( .A(
        my_filter_q_reg_coeff[129]), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_n110) );
  INV_X1 my_filter_adder_mult_0_multiplication_mult_21_U216 ( .A(
        my_filter_q_reg_coeff[130]), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_n109) );
  INV_X1 my_filter_adder_mult_0_multiplication_mult_21_U215 ( .A(
        my_filter_q_reg_coeff[131]), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_n108) );
  INV_X1 my_filter_adder_mult_0_multiplication_mult_21_U214 ( .A(
        my_filter_q_reg_chain_1__7_), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_n92) );
  INV_X1 my_filter_adder_mult_0_multiplication_mult_21_U213 ( .A(
        my_filter_q_reg_chain_1__6_), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_n93) );
  INV_X1 my_filter_adder_mult_0_multiplication_mult_21_U212 ( .A(
        my_filter_q_reg_chain_1__5_), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_n94) );
  INV_X1 my_filter_adder_mult_0_multiplication_mult_21_U211 ( .A(
        my_filter_q_reg_chain_1__4_), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_n95) );
  INV_X1 my_filter_adder_mult_0_multiplication_mult_21_U210 ( .A(
        my_filter_q_reg_chain_1__2_), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_n97) );
  INV_X1 my_filter_adder_mult_0_multiplication_mult_21_U209 ( .A(
        my_filter_q_reg_chain_1__3_), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_n96) );
  AND2_X1 my_filter_adder_mult_0_multiplication_mult_21_U208 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_13__12_), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_13__13_), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_n3) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U207 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n100), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_13__13_) );
  AND2_X1 my_filter_adder_mult_0_multiplication_mult_21_U206 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_13__9_), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_13__10_), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_n50) );
  AND2_X1 my_filter_adder_mult_0_multiplication_mult_21_U205 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_13__7_), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_13__8_), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_n49) );
  AND2_X1 my_filter_adder_mult_0_multiplication_mult_21_U204 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_13__10_), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_13__11_), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_n46) );
  AND2_X1 my_filter_adder_mult_0_multiplication_mult_21_U203 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_13__8_), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_13__9_), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_n47) );
  AND2_X1 my_filter_adder_mult_0_multiplication_mult_21_U202 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_13__6_), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_13__7_), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_n39) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U201 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_12__11_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U200 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_12__10_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U199 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_11__11_) );
  AND2_X1 my_filter_adder_mult_0_multiplication_mult_21_U198 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_13__11_), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_13__12_), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_n52) );
  AND2_X1 my_filter_adder_mult_0_multiplication_mult_21_U197 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_13__5_), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_13__6_), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_n42) );
  AND2_X1 my_filter_adder_mult_0_multiplication_mult_21_U196 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_13__3_), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_13__4_), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_n41) );
  AND2_X1 my_filter_adder_mult_0_multiplication_mult_21_U195 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_13__1_), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_13__2_), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_n40) );
  AND2_X1 my_filter_adder_mult_0_multiplication_mult_21_U194 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_13__4_), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_13__5_), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_n38) );
  AND2_X1 my_filter_adder_mult_0_multiplication_mult_21_U193 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_13__2_), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_13__3_), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_n37) );
  AND2_X1 my_filter_adder_mult_0_multiplication_mult_21_U192 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_13__0_), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_13__1_), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_n36) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U191 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_12__1_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U190 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_10__0_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U189 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_11__0_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U188 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_11__1_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U187 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_10__1_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U186 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_8__0_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U185 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n113), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_9__0_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U184 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n112), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_9__1_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U183 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n110), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_9__3_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U182 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_8__1_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U181 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_8__3_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U180 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_6__0_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U179 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_7__0_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U178 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_7__1_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U177 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_7__3_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U176 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_7__4_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U175 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_7__5_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U174 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_6__1_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U173 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_6__3_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U172 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_6__5_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U171 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_4__0_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U170 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_5__0_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U169 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_5__1_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U168 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_5__3_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U167 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_5__4_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U166 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_5__5_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U165 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_5__6_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U164 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_5__7_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U163 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_4__1_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U162 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_4__3_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U161 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_4__5_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U160 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_2__0_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U159 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_3__0_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U158 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_3__1_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U157 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_3__3_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U156 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_3__4_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U155 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_3__5_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U154 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_3__6_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U153 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_3__7_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U152 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_3__8_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U151 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_3__9_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U150 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_12__9_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U149 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_11__10_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U148 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_12__7_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U147 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_12__8_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U146 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_10__11_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U145 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_11__8_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U144 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_11__9_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U143 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_12__5_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U142 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_12__6_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U141 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_10__9_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U140 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_10__10_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U139 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_11__6_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U138 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_11__7_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U137 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n103), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_9__10_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U136 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n102), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_9__11_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U135 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_12__3_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U134 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_12__4_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U133 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_10__7_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U132 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_10__8_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U131 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_8__11_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U130 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_12__2_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U129 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_11__4_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U128 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_11__5_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U127 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n105), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_9__8_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U126 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n104), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_9__9_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U125 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_11__3_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U124 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_10__5_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U123 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_10__6_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U122 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_8__9_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U121 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_8__10_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U120 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_10__4_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U119 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_11__2_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U118 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n107), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_9__6_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U117 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n106), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_9__7_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U116 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_7__10_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U115 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_7__11_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U114 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n108), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_9__5_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U113 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_10__2_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U112 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_10__3_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U111 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_8__7_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U110 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_8__8_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U109 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_6__11_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U108 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_8__6_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U107 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n111), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_9__2_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U106 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n109), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_9__4_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U105 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_7__8_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U104 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_7__9_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U103 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_7__7_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U102 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_8__2_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U101 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_8__4_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U100 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_8__5_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U99 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_6__9_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U98 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_6__10_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U97 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_6__8_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U96 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_7__2_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U95 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_7__6_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U94 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_5__10_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U93 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_5__11_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U92 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_5__9_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U91 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_6__2_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U90 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_6__4_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U89 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_6__6_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U88 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_6__7_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U87 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_4__11_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U86 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_4__10_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U85 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_5__2_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U84 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_5__8_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U83 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_3__11_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U82 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_4__2_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U81 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_4__4_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U80 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_4__6_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U79 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_4__7_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U78 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_4__8_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U77 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_4__9_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U76 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_3__2_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U75 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_3__10_) );
  AND2_X1 my_filter_adder_mult_0_multiplication_mult_21_U74 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_ab_0__2_), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_ab_1__1_), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_n14) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U73 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_2__1_) );
  AND2_X1 my_filter_adder_mult_0_multiplication_mult_21_U72 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_ab_0__3_), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_ab_1__2_), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_n13) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U71 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_2__2_) );
  AND2_X1 my_filter_adder_mult_0_multiplication_mult_21_U70 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_ab_0__4_), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_ab_1__3_), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_n12) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U69 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_2__3_) );
  AND2_X1 my_filter_adder_mult_0_multiplication_mult_21_U68 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_ab_0__5_), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_ab_1__4_), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_n11) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U67 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_2__4_) );
  AND2_X1 my_filter_adder_mult_0_multiplication_mult_21_U66 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_ab_0__6_), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_ab_1__5_), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_n10) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U65 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_2__5_) );
  AND2_X1 my_filter_adder_mult_0_multiplication_mult_21_U64 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_ab_0__7_), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_ab_1__6_), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_n9) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U63 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_2__6_) );
  AND2_X1 my_filter_adder_mult_0_multiplication_mult_21_U62 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_ab_0__8_), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_ab_1__7_), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_n8) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U61 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_2__7_) );
  AND2_X1 my_filter_adder_mult_0_multiplication_mult_21_U60 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_ab_0__9_), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_ab_1__8_), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_n7) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U59 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_2__8_) );
  AND2_X1 my_filter_adder_mult_0_multiplication_mult_21_U58 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_ab_0__10_), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_ab_1__9_), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_n6) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U57 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_2__9_) );
  AND2_X1 my_filter_adder_mult_0_multiplication_mult_21_U56 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_ab_0__11_), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_ab_1__10_), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_n5) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U55 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_2__10_) );
  AND2_X1 my_filter_adder_mult_0_multiplication_mult_21_U54 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_ab_0__12_), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_ab_1__11_), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_n4) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U52 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_2__11_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U50 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_1__12_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U49 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_1__2_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U47 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_1__3_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U46 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_1__4_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U42 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_1__5_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U41 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_1__6_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U40 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_1__7_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U39 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_1__8_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U38 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_1__9_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U37 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_1__10_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U36 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_1__11_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U14 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_0__2_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U13 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_0__3_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U12 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_0__4_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U11 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_0__5_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U10 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_0__6_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U9 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_0__7_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U8 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_0__8_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U7 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_0__9_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U6 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_0__10_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U5 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_0__11_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U4 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_0__12_) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U3 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n98), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n112), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_ab_1__1_) );
  INV_X1 my_filter_adder_mult_0_multiplication_mult_21_U2 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_13__13_), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_n85) );
  XOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U51 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_13__12_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_13__13_), .Z(
        my_filter_adder_mult_0_multiplication_mult_21_n51) );
  XOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U48 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_13__10_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_13__11_), .Z(
        my_filter_adder_mult_0_multiplication_mult_21_n48) );
  XOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U45 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_13__11_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_13__12_), .Z(
        my_filter_adder_mult_0_multiplication_mult_21_n45) );
  XOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U44 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_13__8_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_13__9_), .Z(
        my_filter_adder_mult_0_multiplication_mult_21_n44) );
  XOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U43 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_13__9_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_13__10_), .Z(
        my_filter_adder_mult_0_multiplication_mult_21_n43) );
  XOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U35 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_13__7_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_13__8_), .Z(
        my_filter_adder_mult_0_multiplication_mult_21_n35) );
  XOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U34 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_13__5_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_13__6_), .Z(
        my_filter_adder_mult_0_multiplication_mult_21_n34) );
  XOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U33 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_13__3_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_13__4_), .Z(
        my_filter_adder_mult_0_multiplication_mult_21_n33) );
  XOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U32 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_13__1_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_13__2_), .Z(
        my_filter_adder_mult_0_multiplication_mult_21_n32) );
  XOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U31 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_13__6_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_13__7_), .Z(
        my_filter_adder_mult_0_multiplication_mult_21_n31) );
  XOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U30 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_13__4_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_13__5_), .Z(
        my_filter_adder_mult_0_multiplication_mult_21_n30) );
  XOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U29 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_13__2_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_13__3_), .Z(
        my_filter_adder_mult_0_multiplication_mult_21_n29) );
  XOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U28 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_13__0_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_13__1_), .Z(
        my_filter_adder_mult_0_multiplication_mult_21_n28) );
  XOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U26 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_1__1_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_ab_0__2_), .Z(
        my_filter_adder_mult_0_multiplication_mult_21_n27) );
  XOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U25 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_1__12_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_ab_0__13_), .Z(
        my_filter_adder_mult_0_multiplication_mult_21_n26) );
  XOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U24 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_1__2_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_ab_0__3_), .Z(
        my_filter_adder_mult_0_multiplication_mult_21_n25) );
  XOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U23 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_1__3_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_ab_0__4_), .Z(
        my_filter_adder_mult_0_multiplication_mult_21_n24) );
  XOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U22 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_1__4_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_ab_0__5_), .Z(
        my_filter_adder_mult_0_multiplication_mult_21_n23) );
  XOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U21 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_1__5_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_ab_0__6_), .Z(
        my_filter_adder_mult_0_multiplication_mult_21_n22) );
  XOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U20 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_1__6_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_ab_0__7_), .Z(
        my_filter_adder_mult_0_multiplication_mult_21_n21) );
  XOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U19 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_1__7_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_ab_0__8_), .Z(
        my_filter_adder_mult_0_multiplication_mult_21_n20) );
  XOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U18 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_1__8_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_ab_0__9_), .Z(
        my_filter_adder_mult_0_multiplication_mult_21_n19) );
  XOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U17 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_1__9_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_ab_0__10_), .Z(
        my_filter_adder_mult_0_multiplication_mult_21_n18) );
  XOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U16 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_1__10_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_ab_0__11_), .Z(
        my_filter_adder_mult_0_multiplication_mult_21_n17) );
  XOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_U15 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_1__11_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_ab_0__12_), .Z(
        my_filter_adder_mult_0_multiplication_mult_21_n16) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S3_2_12 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_2__12_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_n15), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_ab_1__13_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_2__12_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_2__12_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_2_11 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_2__11_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_n4), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_n26), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_2__11_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_2__11_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_2_10 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_2__10_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_n5), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_n16), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_2__10_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_2__10_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_2_9 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_2__9_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_n6), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_n17), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_2__9_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_2__9_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_2_8 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_2__8_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_n7), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_n18), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_2__8_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_2__8_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_2_7 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_2__7_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_n8), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_n19), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_2__7_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_2__7_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_2_6 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_2__6_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_n9), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_n20), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_2__6_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_2__6_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_2_5 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_2__5_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_n10), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_n21), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_2__5_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_2__5_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_2_4 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_2__4_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_n11), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_n22), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_2__4_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_2__4_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_2_3 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_2__3_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_n12), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_n23), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_2__3_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_2__3_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_2_2 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_2__2_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_n13), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_n24), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_2__2_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_2__2_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_2_1 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_2__1_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_n14), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_n25), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_2__1_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_2__1_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S1_2_0 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_2__0_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_1__0_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_n27), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_2__0_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_A1_0_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S3_3_12 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_3__12_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_2__12_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_ab_2__13_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_3__12_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_3__12_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_3_11 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_3__11_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_2__11_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_2__12_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_3__11_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_3__11_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_3_10 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_3__10_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_2__10_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_2__11_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_3__10_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_3__10_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_3_9 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_3__9_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_2__9_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_2__10_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_3__9_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_3__9_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_3_8 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_3__8_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_2__8_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_2__9_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_3__8_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_3__8_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_3_7 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_3__7_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_2__7_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_2__8_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_3__7_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_3__7_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_3_6 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_3__6_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_2__6_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_2__7_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_3__6_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_3__6_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_3_5 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_3__5_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_2__5_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_2__6_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_3__5_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_3__5_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_3_4 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_3__4_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_2__4_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_2__5_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_3__4_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_3__4_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_3_3 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_3__3_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_2__3_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_2__4_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_3__3_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_3__3_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_3_2 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_3__2_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_2__2_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_2__3_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_3__2_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_3__2_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_3_1 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_3__1_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_2__1_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_2__2_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_3__1_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_3__1_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S1_3_0 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_3__0_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_2__0_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_2__1_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_3__0_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_A1_1_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S3_4_12 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_4__12_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_3__12_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_ab_3__13_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_4__12_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_4__12_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_4_11 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_4__11_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_3__11_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_3__12_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_4__11_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_4__11_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_4_10 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_4__10_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_3__10_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_3__11_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_4__10_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_4__10_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_4_9 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_4__9_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_3__9_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_3__10_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_4__9_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_4__9_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_4_8 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_4__8_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_3__8_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_3__9_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_4__8_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_4__8_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_4_7 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_4__7_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_3__7_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_3__8_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_4__7_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_4__7_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_4_6 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_4__6_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_3__6_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_3__7_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_4__6_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_4__6_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_4_5 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_4__5_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_3__5_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_3__6_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_4__5_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_4__5_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_4_4 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_4__4_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_3__4_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_3__5_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_4__4_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_4__4_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_4_3 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_4__3_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_3__3_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_3__4_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_4__3_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_4__3_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_4_2 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_4__2_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_3__2_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_3__3_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_4__2_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_4__2_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_4_1 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_4__1_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_3__1_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_3__2_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_4__1_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_4__1_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S1_4_0 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_4__0_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_3__0_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_3__1_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_4__0_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_A1_2_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S3_5_12 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_5__12_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_4__12_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_ab_4__13_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_5__12_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_5__12_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_5_11 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_5__11_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_4__11_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_4__12_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_5__11_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_5__11_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_5_10 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_5__10_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_4__10_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_4__11_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_5__10_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_5__10_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_5_9 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_5__9_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_4__9_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_4__10_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_5__9_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_5__9_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_5_8 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_5__8_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_4__8_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_4__9_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_5__8_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_5__8_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_5_7 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_5__7_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_4__7_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_4__8_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_5__7_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_5__7_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_5_6 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_5__6_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_4__6_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_4__7_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_5__6_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_5__6_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_5_5 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_5__5_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_4__5_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_4__6_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_5__5_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_5__5_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_5_4 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_5__4_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_4__4_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_4__5_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_5__4_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_5__4_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_5_3 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_5__3_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_4__3_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_4__4_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_5__3_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_5__3_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_5_2 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_5__2_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_4__2_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_4__3_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_5__2_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_5__2_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_5_1 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_5__1_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_4__1_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_4__2_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_5__1_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_5__1_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S1_5_0 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_5__0_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_4__0_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_4__1_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_5__0_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_A1_3_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S3_6_12 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_6__12_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_5__12_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_ab_5__13_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_6__12_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_6__12_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_6_11 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_6__11_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_5__11_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_5__12_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_6__11_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_6__11_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_6_10 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_6__10_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_5__10_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_5__11_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_6__10_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_6__10_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_6_9 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_6__9_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_5__9_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_5__10_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_6__9_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_6__9_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_6_8 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_6__8_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_5__8_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_5__9_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_6__8_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_6__8_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_6_7 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_6__7_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_5__7_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_5__8_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_6__7_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_6__7_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_6_6 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_6__6_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_5__6_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_5__7_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_6__6_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_6__6_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_6_5 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_6__5_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_5__5_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_5__6_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_6__5_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_6__5_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_6_4 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_6__4_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_5__4_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_5__5_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_6__4_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_6__4_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_6_3 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_6__3_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_5__3_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_5__4_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_6__3_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_6__3_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_6_2 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_6__2_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_5__2_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_5__3_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_6__2_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_6__2_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_6_1 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_6__1_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_5__1_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_5__2_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_6__1_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_6__1_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S1_6_0 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_6__0_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_5__0_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_5__1_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_6__0_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_A1_4_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S3_7_12 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_7__12_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_6__12_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_ab_6__13_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_7__12_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_7__12_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_7_11 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_7__11_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_6__11_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_6__12_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_7__11_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_7__11_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_7_10 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_7__10_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_6__10_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_6__11_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_7__10_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_7__10_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_7_9 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_7__9_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_6__9_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_6__10_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_7__9_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_7__9_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_7_8 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_7__8_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_6__8_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_6__9_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_7__8_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_7__8_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_7_7 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_7__7_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_6__7_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_6__8_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_7__7_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_7__7_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_7_6 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_7__6_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_6__6_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_6__7_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_7__6_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_7__6_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_7_5 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_7__5_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_6__5_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_6__6_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_7__5_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_7__5_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_7_4 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_7__4_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_6__4_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_6__5_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_7__4_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_7__4_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_7_3 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_7__3_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_6__3_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_6__4_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_7__3_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_7__3_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_7_2 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_7__2_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_6__2_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_6__3_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_7__2_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_7__2_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_7_1 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_7__1_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_6__1_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_6__2_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_7__1_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_7__1_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S1_7_0 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_7__0_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_6__0_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_6__1_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_7__0_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_A1_5_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S3_8_12 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_8__12_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_7__12_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_ab_7__13_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_8__12_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_8__12_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_8_11 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_8__11_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_7__11_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_7__12_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_8__11_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_8__11_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_8_10 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_8__10_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_7__10_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_7__11_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_8__10_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_8__10_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_8_9 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_8__9_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_7__9_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_7__10_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_8__9_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_8__9_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_8_8 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_8__8_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_7__8_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_7__9_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_8__8_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_8__8_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_8_7 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_8__7_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_7__7_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_7__8_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_8__7_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_8__7_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_8_6 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_8__6_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_7__6_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_7__7_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_8__6_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_8__6_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_8_5 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_8__5_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_7__5_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_7__6_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_8__5_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_8__5_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_8_4 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_8__4_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_7__4_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_7__5_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_8__4_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_8__4_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_8_3 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_8__3_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_7__3_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_7__4_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_8__3_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_8__3_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_8_2 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_8__2_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_7__2_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_7__3_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_8__2_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_8__2_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_8_1 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_8__1_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_7__1_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_7__2_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_8__1_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_8__1_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S1_8_0 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_8__0_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_7__0_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_7__1_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_8__0_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_A1_6_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S3_9_12 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_9__12_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_8__12_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_ab_8__13_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_9__12_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_9__12_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_9_11 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_9__11_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_8__11_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_8__12_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_9__11_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_9__11_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_9_10 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_9__10_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_8__10_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_8__11_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_9__10_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_9__10_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_9_9 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_9__9_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_8__9_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_8__10_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_9__9_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_9__9_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_9_8 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_9__8_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_8__8_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_8__9_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_9__8_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_9__8_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_9_7 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_9__7_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_8__7_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_8__8_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_9__7_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_9__7_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_9_6 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_9__6_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_8__6_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_8__7_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_9__6_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_9__6_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_9_5 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_9__5_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_8__5_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_8__6_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_9__5_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_9__5_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_9_4 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_9__4_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_8__4_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_8__5_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_9__4_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_9__4_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_9_3 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_9__3_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_8__3_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_8__4_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_9__3_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_9__3_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_9_2 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_9__2_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_8__2_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_8__3_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_9__2_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_9__2_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_9_1 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_9__1_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_8__1_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_8__2_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_9__1_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_9__1_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S1_9_0 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_9__0_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_8__0_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_8__1_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_9__0_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_A1_7_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S3_10_12 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_10__12_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_9__12_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_ab_9__13_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_10__12_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_10__12_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_10_11 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_10__11_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_9__11_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_9__12_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_10__11_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_10__11_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_10_10 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_10__10_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_9__10_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_9__11_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_10__10_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_10__10_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_10_9 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_10__9_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_9__9_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_9__10_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_10__9_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_10__9_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_10_8 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_10__8_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_9__8_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_9__9_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_10__8_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_10__8_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_10_7 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_10__7_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_9__7_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_9__8_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_10__7_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_10__7_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_10_6 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_10__6_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_9__6_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_9__7_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_10__6_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_10__6_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_10_5 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_10__5_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_9__5_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_9__6_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_10__5_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_10__5_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_10_4 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_10__4_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_9__4_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_9__5_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_10__4_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_10__4_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_10_3 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_10__3_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_9__3_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_9__4_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_10__3_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_10__3_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_10_2 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_10__2_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_9__2_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_9__3_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_10__2_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_10__2_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_10_1 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_10__1_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_9__1_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_9__2_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_10__1_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_10__1_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S1_10_0 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_10__0_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_9__0_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_9__1_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_10__0_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_A1_8_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S3_11_12 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_11__12_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_10__12_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_ab_10__13_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_11__12_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_11__12_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_11_11 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_11__11_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_10__11_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_10__12_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_11__11_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_11__11_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_11_10 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_11__10_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_10__10_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_10__11_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_11__10_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_11__10_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_11_9 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_11__9_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_10__9_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_10__10_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_11__9_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_11__9_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_11_8 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_11__8_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_10__8_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_10__9_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_11__8_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_11__8_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_11_7 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_11__7_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_10__7_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_10__8_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_11__7_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_11__7_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_11_6 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_11__6_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_10__6_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_10__7_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_11__6_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_11__6_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_11_5 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_11__5_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_10__5_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_10__6_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_11__5_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_11__5_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_11_4 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_11__4_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_10__4_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_10__5_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_11__4_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_11__4_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_11_3 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_11__3_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_10__3_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_10__4_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_11__3_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_11__3_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_11_2 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_11__2_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_10__2_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_10__3_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_11__2_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_11__2_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_11_1 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_11__1_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_10__1_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_10__2_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_11__1_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_11__1_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S1_11_0 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_11__0_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_10__0_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_10__1_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_11__0_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_A1_9_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S3_12_12 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_12__12_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_11__12_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_ab_11__13_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_12__12_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_12__12_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_12_11 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_12__11_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_11__11_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_11__12_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_12__11_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_12__11_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_12_10 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_12__10_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_11__10_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_11__11_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_12__10_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_12__10_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_12_9 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_12__9_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_11__9_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_11__10_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_12__9_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_12__9_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_12_8 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_12__8_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_11__8_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_11__9_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_12__8_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_12__8_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_12_7 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_12__7_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_11__7_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_11__8_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_12__7_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_12__7_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_12_6 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_12__6_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_11__6_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_11__7_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_12__6_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_12__6_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_12_5 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_12__5_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_11__5_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_11__6_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_12__5_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_12__5_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_12_4 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_12__4_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_11__4_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_11__5_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_12__4_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_12__4_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_12_3 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_12__3_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_11__3_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_11__4_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_12__3_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_12__3_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_12_2 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_12__2_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_11__2_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_11__3_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_12__2_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_12__2_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S2_12_1 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_12__1_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_11__1_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_11__2_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_12__1_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_12__1_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S1_12_0 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_12__0_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_11__0_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_11__1_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_12__0_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_A1_10_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S14_13 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_n86), .B(
        my_filter_adder_mult_0_multiplication_mult_21_n100), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_ab_13__13_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_13__13_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_13__13_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S5_12 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_13__12_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_12__12_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_ab_12__13_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_13__12_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_13__12_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S4_11 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_13__11_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_12__11_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_12__12_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_13__11_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_13__11_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S4_10 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_13__10_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_12__10_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_12__11_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_13__10_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_13__10_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S4_9 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_13__9_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_12__9_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_12__10_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_13__9_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_13__9_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S4_8 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_13__8_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_12__8_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_12__9_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_13__8_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_13__8_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S4_7 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_13__7_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_12__7_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_12__8_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_13__7_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_13__7_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S4_6 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_13__6_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_12__6_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_12__7_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_13__6_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_13__6_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S4_5 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_13__5_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_12__5_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_12__6_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_13__5_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_13__5_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S4_4 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_13__4_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_12__4_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_12__5_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_13__4_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_13__4_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S4_3 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_13__3_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_12__3_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_12__4_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_13__3_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_13__3_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S4_2 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_13__2_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_12__2_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_12__3_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_13__2_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_13__2_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S4_1 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_13__1_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_12__1_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_12__2_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_13__1_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_13__1_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S4_0 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_ab_13__0_), .B(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_12__0_), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_12__1_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_CARRYB_13__0_), .S(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_13__0_) );
  FA_X1 my_filter_adder_mult_0_multiplication_mult_21_S14_13_0 ( .A(
        my_filter_q_reg_chain_1__13_), .B(my_filter_q_reg_coeff[139]), .CI(
        my_filter_adder_mult_0_multiplication_mult_21_SUMB_13__0_), .CO(
        my_filter_adder_mult_0_multiplication_mult_21_A2_12_), .S(
        my_filter_adder_mult_0_res_mult[0]) );
  NAND2_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U72 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_A2_12_), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n28), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n56) );
  INV_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U71 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n59), .ZN(
        my_filter_adder_mult_0_res_mult[1]) );
  OAI21_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U70 ( .B1(
        my_filter_adder_mult_0_multiplication_mult_21_A2_12_), .B2(
        my_filter_adder_mult_0_multiplication_mult_21_n28), .A(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n56), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n59) );
  AND2_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U69 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n50), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n48), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n20) );
  AND2_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U68 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n49), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n44), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n28) );
  NAND2_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U66 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n46), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n45), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n17) );
  NAND2_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U65 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n47), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n43), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n25) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U64 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n46), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n45), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n15) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U63 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n47), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n43), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n23) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U61 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n50), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n48), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n21) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U60 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n49), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n44), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n29) );
  AND2_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U59 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n42), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n31), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n36) );
  AND2_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U58 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n41), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n30), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n44) );
  AND2_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U56 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n40), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n29), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n52) );
  NAND2_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U55 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n39), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n35), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n33) );
  NAND2_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U54 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n38), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n34), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n41) );
  NAND2_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U53 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n37), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n33), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n49) );
  NAND2_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U51 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n36), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n32), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n57) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U50 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n39), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n35), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n31) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U49 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n38), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n34), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n39) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U48 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n37), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n33), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n47) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U46 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n36), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n32), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n55) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U45 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n42), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n31), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n37) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U44 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n41), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n30), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n45) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U43 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_n40), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_n29), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n53) );
  OAI21_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U41 ( .B1(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n55), .B2(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n56), .A(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n57), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n51) );
  INV_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U40 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n15), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n62) );
  INV_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U39 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n23), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n64) );
  INV_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U38 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n31), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n70) );
  INV_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U36 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n39), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n68) );
  NAND2_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U35 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n68), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n41), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n42) );
  INV_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U34 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n47), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n66) );
  NAND2_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U33 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n66), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n49), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n50) );
  INV_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U31 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n55), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n60) );
  NAND2_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U30 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n60), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n57), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n58) );
  NAND2_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U29 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n62), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n17), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n18) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U28 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n20), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n21), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n22) );
  NAND2_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U26 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n64), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n25), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n26) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U25 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n28), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n29), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n30) );
  NAND2_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U24 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n70), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n33), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n34) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U23 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n36), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n37), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n38) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U21 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n44), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n45), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n46) );
  NOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U20 ( .A1(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n52), .A2(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n53), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n54) );
  OAI21_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U19 ( .B1(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n15), .B2(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n16), .A(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n17), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n13) );
  OAI21_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U18 ( .B1(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n23), .B2(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n24), .A(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n25), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n19) );
  OAI21_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U16 ( .B1(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n31), .B2(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n32), .A(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n33), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n27) );
  OAI21_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U13 ( .B1(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n39), .B2(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n40), .A(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n41), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n35) );
  OAI21_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U12 ( .B1(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n47), .B2(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n48), .A(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n49), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n43) );
  INV_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U11 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n21), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n63) );
  AOI21_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U10 ( .B1(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n63), .B2(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n19), .A(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n20), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n16) );
  INV_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U9 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n29), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n71) );
  AOI21_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U8 ( .B1(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n71), .B2(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n27), .A(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n28), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n24) );
  INV_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U7 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n37), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n69) );
  AOI21_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U6 ( .B1(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n69), .B2(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n35), .A(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n36), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n32) );
  INV_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U5 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n45), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n67) );
  AOI21_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U4 ( .B1(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n67), .B2(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n43), .A(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n44), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n40) );
  INV_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U3 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n53), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n65) );
  AOI21_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U2 ( .B1(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n65), .B2(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n51), .A(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n52), .ZN(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n48) );
  XOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U67 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n56), .B(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n58), .Z(
        my_filter_adder_mult_0_res_mult[2]) );
  XOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U62 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n51), .B(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n54), .Z(
        my_filter_adder_mult_0_res_mult[3]) );
  XOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U57 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n50), .B(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n48), .Z(
        my_filter_adder_mult_0_res_mult[4]) );
  XOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U52 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n43), .B(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n46), .Z(
        my_filter_adder_mult_0_res_mult[5]) );
  XOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U47 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n42), .B(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n40), .Z(
        my_filter_adder_mult_0_res_mult[6]) );
  XOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U42 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n35), .B(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n38), .Z(
        my_filter_adder_mult_0_res_mult[7]) );
  XOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U37 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n34), .B(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n32), .Z(
        my_filter_adder_mult_0_res_mult[8]) );
  XOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U32 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n27), .B(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n30), .Z(
        my_filter_adder_mult_0_res_mult[9]) );
  XOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U27 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n26), .B(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n24), .Z(
        my_filter_adder_mult_0_res_mult[10]) );
  XOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U22 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n19), .B(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n22), .Z(
        my_filter_adder_mult_0_res_mult[11]) );
  XOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U17 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n18), .B(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n16), .Z(
        my_filter_adder_mult_0_res_mult[12]) );
  XOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U15 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_n52), .B(
        my_filter_adder_mult_0_multiplication_mult_21_n51), .Z(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n14) );
  XOR2_X1 my_filter_adder_mult_0_multiplication_mult_21_FS_1_U14 ( .A(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n13), .B(
        my_filter_adder_mult_0_multiplication_mult_21_FS_1_n14), .Z(
        my_filter_adder_mult_0_res_mult[13]) );
  AND2_X1 my_filter_adder_mult_0_addition_add_19_U1 ( .A1(
        my_filter_data_sum[140]), .A2(my_filter_adder_mult_0_res_mult[0]), 
        .ZN(my_filter_adder_mult_0_addition_add_19_n1) );
  XOR2_X1 my_filter_adder_mult_0_addition_add_19_U2 ( .A(
        my_filter_data_sum[140]), .B(my_filter_adder_mult_0_res_mult[0]), .Z(
        my_filter_data_sum[126]) );
  FA_X1 my_filter_adder_mult_0_addition_add_19_U1_1 ( .A(
        my_filter_adder_mult_0_res_mult[1]), .B(my_filter_data_sum[141]), .CI(
        my_filter_adder_mult_0_addition_add_19_n1), .CO(
        my_filter_adder_mult_0_addition_add_19_carry[2]), .S(
        my_filter_data_sum[127]) );
  FA_X1 my_filter_adder_mult_0_addition_add_19_U1_2 ( .A(
        my_filter_adder_mult_0_res_mult[2]), .B(my_filter_data_sum[142]), .CI(
        my_filter_adder_mult_0_addition_add_19_carry[2]), .CO(
        my_filter_adder_mult_0_addition_add_19_carry[3]), .S(
        my_filter_data_sum[128]) );
  FA_X1 my_filter_adder_mult_0_addition_add_19_U1_3 ( .A(
        my_filter_adder_mult_0_res_mult[3]), .B(my_filter_data_sum[143]), .CI(
        my_filter_adder_mult_0_addition_add_19_carry[3]), .CO(
        my_filter_adder_mult_0_addition_add_19_carry[4]), .S(
        my_filter_data_sum[129]) );
  FA_X1 my_filter_adder_mult_0_addition_add_19_U1_4 ( .A(
        my_filter_adder_mult_0_res_mult[4]), .B(my_filter_data_sum[144]), .CI(
        my_filter_adder_mult_0_addition_add_19_carry[4]), .CO(
        my_filter_adder_mult_0_addition_add_19_carry[5]), .S(
        my_filter_data_sum[130]) );
  FA_X1 my_filter_adder_mult_0_addition_add_19_U1_5 ( .A(
        my_filter_adder_mult_0_res_mult[5]), .B(my_filter_data_sum[145]), .CI(
        my_filter_adder_mult_0_addition_add_19_carry[5]), .CO(
        my_filter_adder_mult_0_addition_add_19_carry[6]), .S(
        my_filter_data_sum[131]) );
  FA_X1 my_filter_adder_mult_0_addition_add_19_U1_6 ( .A(
        my_filter_adder_mult_0_res_mult[6]), .B(my_filter_data_sum[146]), .CI(
        my_filter_adder_mult_0_addition_add_19_carry[6]), .CO(
        my_filter_adder_mult_0_addition_add_19_carry[7]), .S(
        my_filter_data_sum[132]) );
  FA_X1 my_filter_adder_mult_0_addition_add_19_U1_7 ( .A(
        my_filter_adder_mult_0_res_mult[7]), .B(my_filter_data_sum[147]), .CI(
        my_filter_adder_mult_0_addition_add_19_carry[7]), .CO(
        my_filter_adder_mult_0_addition_add_19_carry[8]), .S(
        my_filter_data_sum[133]) );
  FA_X1 my_filter_adder_mult_0_addition_add_19_U1_8 ( .A(
        my_filter_adder_mult_0_res_mult[8]), .B(my_filter_data_sum[148]), .CI(
        my_filter_adder_mult_0_addition_add_19_carry[8]), .CO(
        my_filter_adder_mult_0_addition_add_19_carry[9]), .S(
        my_filter_data_sum[134]) );
  FA_X1 my_filter_adder_mult_0_addition_add_19_U1_9 ( .A(
        my_filter_adder_mult_0_res_mult[9]), .B(my_filter_data_sum[149]), .CI(
        my_filter_adder_mult_0_addition_add_19_carry[9]), .CO(
        my_filter_adder_mult_0_addition_add_19_carry[10]), .S(
        my_filter_data_sum[135]) );
  FA_X1 my_filter_adder_mult_0_addition_add_19_U1_10 ( .A(
        my_filter_adder_mult_0_res_mult[10]), .B(my_filter_data_sum[150]), 
        .CI(my_filter_adder_mult_0_addition_add_19_carry[10]), .CO(
        my_filter_adder_mult_0_addition_add_19_carry[11]), .S(
        my_filter_data_sum[136]) );
  FA_X1 my_filter_adder_mult_0_addition_add_19_U1_11 ( .A(
        my_filter_adder_mult_0_res_mult[11]), .B(my_filter_data_sum[151]), 
        .CI(my_filter_adder_mult_0_addition_add_19_carry[11]), .CO(
        my_filter_adder_mult_0_addition_add_19_carry[12]), .S(
        my_filter_data_sum[137]) );
  FA_X1 my_filter_adder_mult_0_addition_add_19_U1_12 ( .A(
        my_filter_adder_mult_0_res_mult[12]), .B(my_filter_data_sum[152]), 
        .CI(my_filter_adder_mult_0_addition_add_19_carry[12]), .CO(
        my_filter_adder_mult_0_addition_add_19_carry[13]), .S(
        my_filter_data_sum[138]) );
  FA_X1 my_filter_adder_mult_0_addition_add_19_U1_13 ( .A(
        my_filter_adder_mult_0_res_mult[13]), .B(my_filter_data_sum[153]), 
        .CI(my_filter_adder_mult_0_addition_add_19_carry[13]), .S(
        my_filter_data_sum[139]) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U276 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_12__12_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U275 ( .A1(
        my_filter_q_reg_chain_2__11_), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_11__13_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U274 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_11__12_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U273 ( .A1(
        my_filter_q_reg_chain_2__10_), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_10__13_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U272 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_10__12_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U271 ( .A1(
        my_filter_q_reg_chain_2__9_), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_9__13_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U270 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n101), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_9__12_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U269 ( .A1(
        my_filter_q_reg_chain_2__8_), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_8__13_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U268 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_8__12_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U267 ( .A1(
        my_filter_q_reg_chain_2__7_), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_7__13_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U266 ( .A1(
        my_filter_q_reg_coeff[123]), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_13__11_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U265 ( .A1(
        my_filter_q_reg_coeff[122]), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_13__10_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U264 ( .A1(
        my_filter_q_reg_coeff[120]), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_13__8_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U263 ( .A1(
        my_filter_q_reg_coeff[121]), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_13__9_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U262 ( .A1(
        my_filter_q_reg_coeff[119]), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_13__7_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U261 ( .A1(
        my_filter_q_reg_coeff[124]), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_13__12_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U260 ( .A1(
        my_filter_q_reg_chain_2__12_), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_12__13_) );
  INV_X1 my_filter_adder_mult_1_multiplication_mult_21_U259 ( .A(
        my_filter_q_reg_chain_2__9_), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_n90) );
  INV_X1 my_filter_adder_mult_1_multiplication_mult_21_U258 ( .A(
        my_filter_q_reg_chain_2__12_), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_n87) );
  INV_X1 my_filter_adder_mult_1_multiplication_mult_21_U257 ( .A(
        my_filter_q_reg_chain_2__11_), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_n88) );
  INV_X1 my_filter_adder_mult_1_multiplication_mult_21_U256 ( .A(
        my_filter_q_reg_chain_2__10_), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_n89) );
  INV_X1 my_filter_adder_mult_1_multiplication_mult_21_U255 ( .A(
        my_filter_q_reg_chain_2__8_), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_n91) );
  INV_X1 my_filter_adder_mult_1_multiplication_mult_21_U254 ( .A(
        my_filter_q_reg_chain_2__7_), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_n92) );
  INV_X1 my_filter_adder_mult_1_multiplication_mult_21_U253 ( .A(
        my_filter_q_reg_chain_2__13_), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_n86) );
  AND2_X1 my_filter_adder_mult_1_multiplication_mult_21_U252 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_ab_0__13_), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_ab_1__12_), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_n15) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U251 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_2__12_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U250 ( .A1(
        my_filter_q_reg_chain_2__1_), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_1__13_) );
  AND3_X1 my_filter_adder_mult_1_multiplication_mult_21_U249 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_ab_1__1_), .A2(
        my_filter_q_reg_coeff[112]), .A3(my_filter_q_reg_chain_2__0_), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_1__0_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U248 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_12__0_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U247 ( .A1(
        my_filter_q_reg_coeff[112]), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_13__0_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U246 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_7__12_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U245 ( .A1(
        my_filter_q_reg_chain_2__6_), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_6__13_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U244 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_6__12_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U243 ( .A1(
        my_filter_q_reg_chain_2__5_), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_5__13_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U242 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_5__12_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U241 ( .A1(
        my_filter_q_reg_chain_2__4_), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_4__13_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U240 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_4__12_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U239 ( .A1(
        my_filter_q_reg_chain_2__3_), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_3__13_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U238 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_3__12_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U237 ( .A1(
        my_filter_q_reg_chain_2__2_), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_2__13_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U236 ( .A1(
        my_filter_q_reg_coeff[118]), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_13__6_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U235 ( .A1(
        my_filter_q_reg_coeff[116]), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_13__4_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U234 ( .A1(
        my_filter_q_reg_coeff[117]), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_13__5_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U233 ( .A1(
        my_filter_q_reg_coeff[113]), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_13__1_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U232 ( .A1(
        my_filter_q_reg_coeff[114]), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_13__2_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U231 ( .A1(
        my_filter_q_reg_coeff[115]), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_13__3_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U230 ( .A1(
        my_filter_q_reg_chain_2__0_), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_0__13_) );
  INV_X1 my_filter_adder_mult_1_multiplication_mult_21_U229 ( .A(
        my_filter_q_reg_coeff[125]), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_n100) );
  INV_X1 my_filter_adder_mult_1_multiplication_mult_21_U228 ( .A(
        my_filter_q_reg_coeff[112]), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_n113) );
  INV_X1 my_filter_adder_mult_1_multiplication_mult_21_U227 ( .A(
        my_filter_q_reg_chain_2__0_), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_n99) );
  INV_X1 my_filter_adder_mult_1_multiplication_mult_21_U226 ( .A(
        my_filter_q_reg_coeff[113]), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_n112) );
  INV_X1 my_filter_adder_mult_1_multiplication_mult_21_U225 ( .A(
        my_filter_q_reg_chain_2__1_), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_n98) );
  INV_X1 my_filter_adder_mult_1_multiplication_mult_21_U224 ( .A(
        my_filter_q_reg_coeff[124]), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_n101) );
  INV_X1 my_filter_adder_mult_1_multiplication_mult_21_U223 ( .A(
        my_filter_q_reg_coeff[122]), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_n103) );
  INV_X1 my_filter_adder_mult_1_multiplication_mult_21_U222 ( .A(
        my_filter_q_reg_coeff[123]), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_n102) );
  INV_X1 my_filter_adder_mult_1_multiplication_mult_21_U221 ( .A(
        my_filter_q_reg_coeff[120]), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_n105) );
  INV_X1 my_filter_adder_mult_1_multiplication_mult_21_U220 ( .A(
        my_filter_q_reg_coeff[121]), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_n104) );
  INV_X1 my_filter_adder_mult_1_multiplication_mult_21_U219 ( .A(
        my_filter_q_reg_coeff[117]), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_n108) );
  INV_X1 my_filter_adder_mult_1_multiplication_mult_21_U218 ( .A(
        my_filter_q_reg_coeff[118]), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_n107) );
  INV_X1 my_filter_adder_mult_1_multiplication_mult_21_U217 ( .A(
        my_filter_q_reg_coeff[119]), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_n106) );
  INV_X1 my_filter_adder_mult_1_multiplication_mult_21_U216 ( .A(
        my_filter_q_reg_coeff[114]), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_n111) );
  INV_X1 my_filter_adder_mult_1_multiplication_mult_21_U215 ( .A(
        my_filter_q_reg_coeff[115]), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_n110) );
  INV_X1 my_filter_adder_mult_1_multiplication_mult_21_U214 ( .A(
        my_filter_q_reg_coeff[116]), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_n109) );
  INV_X1 my_filter_adder_mult_1_multiplication_mult_21_U213 ( .A(
        my_filter_q_reg_chain_2__6_), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_n93) );
  INV_X1 my_filter_adder_mult_1_multiplication_mult_21_U212 ( .A(
        my_filter_q_reg_chain_2__5_), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_n94) );
  INV_X1 my_filter_adder_mult_1_multiplication_mult_21_U211 ( .A(
        my_filter_q_reg_chain_2__4_), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_n95) );
  INV_X1 my_filter_adder_mult_1_multiplication_mult_21_U210 ( .A(
        my_filter_q_reg_chain_2__2_), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_n97) );
  INV_X1 my_filter_adder_mult_1_multiplication_mult_21_U209 ( .A(
        my_filter_q_reg_chain_2__3_), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_n96) );
  AND2_X1 my_filter_adder_mult_1_multiplication_mult_21_U208 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_13__12_), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_13__13_), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_n3) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U207 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n100), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_13__13_) );
  AND2_X1 my_filter_adder_mult_1_multiplication_mult_21_U206 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_13__9_), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_13__10_), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_n51) );
  AND2_X1 my_filter_adder_mult_1_multiplication_mult_21_U205 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_13__7_), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_13__8_), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_n50) );
  AND2_X1 my_filter_adder_mult_1_multiplication_mult_21_U204 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_13__5_), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_13__6_), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_n41) );
  AND2_X1 my_filter_adder_mult_1_multiplication_mult_21_U203 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_13__10_), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_13__11_), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_n47) );
  AND2_X1 my_filter_adder_mult_1_multiplication_mult_21_U202 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_13__8_), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_13__9_), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_n46) );
  AND2_X1 my_filter_adder_mult_1_multiplication_mult_21_U201 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_13__6_), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_13__7_), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_n45) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U200 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_12__11_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U199 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_12__9_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U198 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_12__10_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U197 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_11__10_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U196 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_11__11_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U195 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_12__8_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U194 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_10__11_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U193 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_11__9_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U192 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_10__10_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U191 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n102), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_9__11_) );
  AND2_X1 my_filter_adder_mult_1_multiplication_mult_21_U190 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_13__3_), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_13__4_), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_n33) );
  AND2_X1 my_filter_adder_mult_1_multiplication_mult_21_U189 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_13__1_), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_13__2_), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_n40) );
  AND2_X1 my_filter_adder_mult_1_multiplication_mult_21_U188 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_13__4_), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_13__5_), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_n39) );
  AND2_X1 my_filter_adder_mult_1_multiplication_mult_21_U187 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_13__2_), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_13__3_), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_n38) );
  AND2_X1 my_filter_adder_mult_1_multiplication_mult_21_U186 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_13__0_), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_13__1_), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_n37) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U185 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_12__1_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U184 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_10__0_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U183 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_11__0_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U182 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_11__1_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U181 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_10__1_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U180 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_8__0_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U179 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n113), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_9__0_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U178 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n112), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_9__1_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U177 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n110), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_9__3_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U176 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_8__1_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U175 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_8__3_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U174 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_6__0_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U173 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_7__0_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U172 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_7__1_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U171 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_7__3_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U170 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_7__4_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U169 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_7__5_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U168 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_6__1_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U167 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_6__3_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U166 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_6__5_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U165 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_4__0_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U164 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_5__0_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U163 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_5__1_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U162 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_5__3_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U161 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_5__4_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U160 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_5__5_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U159 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_5__6_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U158 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_4__1_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U157 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_4__3_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U156 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_4__5_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U155 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_2__0_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U154 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_3__0_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U153 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_3__1_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U152 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_3__3_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U151 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_3__4_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U150 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_3__5_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U149 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_3__6_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U148 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_3__7_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U147 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_12__7_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U146 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_11__8_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U145 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_12__5_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U144 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_12__6_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U143 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_10__9_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U142 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_11__6_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U141 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_11__7_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U140 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n103), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_9__10_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U139 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_12__2_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U138 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_12__3_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U137 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_12__4_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U136 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_10__7_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U135 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_10__8_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U134 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_8__11_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U133 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_11__3_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U132 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_11__4_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U131 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_11__5_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U130 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n105), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_9__8_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U129 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n104), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_9__9_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U128 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_10__4_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U127 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_10__5_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U126 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_10__6_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U125 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_8__9_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U124 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_8__10_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U123 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_11__2_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U122 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n108), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_9__5_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U121 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n107), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_9__6_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U120 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n106), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_9__7_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U119 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_7__10_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U118 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_7__11_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U117 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_10__2_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U116 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_10__3_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U115 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_8__6_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U114 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_8__7_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U113 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_8__8_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U112 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_6__11_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U111 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n111), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_9__2_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U110 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n109), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_9__4_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U109 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_7__7_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U108 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_7__8_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U107 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_7__9_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U106 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_8__2_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U105 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_8__4_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U104 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_8__5_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U103 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_6__8_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U102 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_6__9_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U101 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_6__10_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U100 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_7__2_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U99 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_7__6_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U98 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_5__9_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U97 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_5__10_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U96 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_5__11_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U95 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_6__2_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U94 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_6__4_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U93 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_6__6_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U92 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_6__7_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U91 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_4__10_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U90 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_4__11_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U89 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_5__2_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U88 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_5__7_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U87 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_5__8_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U86 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_3__11_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U85 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_4__2_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U84 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_4__4_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U83 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_4__6_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U82 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_4__7_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U81 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_4__8_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U80 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_4__9_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U79 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_3__2_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U78 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_3__8_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U77 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_3__9_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U76 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_3__10_) );
  AND2_X1 my_filter_adder_mult_1_multiplication_mult_21_U75 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_ab_0__2_), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_ab_1__1_), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_n14) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U74 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_2__1_) );
  AND2_X1 my_filter_adder_mult_1_multiplication_mult_21_U73 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_ab_0__3_), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_ab_1__2_), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_n13) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U72 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_2__2_) );
  AND2_X1 my_filter_adder_mult_1_multiplication_mult_21_U71 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_ab_0__4_), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_ab_1__3_), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_n12) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U70 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_2__3_) );
  AND2_X1 my_filter_adder_mult_1_multiplication_mult_21_U69 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_ab_0__5_), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_ab_1__4_), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_n11) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U68 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_2__4_) );
  AND2_X1 my_filter_adder_mult_1_multiplication_mult_21_U67 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_ab_0__6_), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_ab_1__5_), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_n10) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U66 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_2__5_) );
  AND2_X1 my_filter_adder_mult_1_multiplication_mult_21_U65 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_ab_0__7_), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_ab_1__6_), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_n9) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U64 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_2__6_) );
  AND2_X1 my_filter_adder_mult_1_multiplication_mult_21_U63 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_ab_0__8_), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_ab_1__7_), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_n8) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U62 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_2__7_) );
  AND2_X1 my_filter_adder_mult_1_multiplication_mult_21_U61 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_ab_0__9_), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_ab_1__8_), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_n7) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U60 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_2__8_) );
  AND2_X1 my_filter_adder_mult_1_multiplication_mult_21_U59 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_ab_0__10_), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_ab_1__9_), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_n6) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U58 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_2__9_) );
  AND2_X1 my_filter_adder_mult_1_multiplication_mult_21_U57 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_ab_0__11_), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_ab_1__10_), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_n5) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U56 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_2__10_) );
  AND2_X1 my_filter_adder_mult_1_multiplication_mult_21_U55 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_ab_0__12_), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_ab_1__11_), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_n4) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U54 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_2__11_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U52 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_1__12_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U51 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_1__2_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U50 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_1__3_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U47 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_1__4_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U46 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_1__5_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U45 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_1__6_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U41 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_1__7_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U40 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_1__8_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U39 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_1__9_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U38 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_1__10_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U37 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_1__11_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U33 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_0__2_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U14 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_0__3_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U13 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_0__4_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U12 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_0__5_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U11 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_0__6_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U10 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_0__7_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U9 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_0__8_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U8 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_0__9_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U7 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_0__10_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U6 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_0__11_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U5 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_0__12_) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U4 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n98), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n112), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_ab_1__1_) );
  AND2_X1 my_filter_adder_mult_1_multiplication_mult_21_U3 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_13__11_), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_13__12_), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_n52) );
  INV_X1 my_filter_adder_mult_1_multiplication_mult_21_U2 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_13__13_), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_n85) );
  XOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U49 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_13__10_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_13__11_), .Z(
        my_filter_adder_mult_1_multiplication_mult_21_n49) );
  XOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U48 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_13__7_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_13__8_), .Z(
        my_filter_adder_mult_1_multiplication_mult_21_n48) );
  XOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U44 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_13__11_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_13__12_), .Z(
        my_filter_adder_mult_1_multiplication_mult_21_n44) );
  XOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U43 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_13__8_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_13__9_), .Z(
        my_filter_adder_mult_1_multiplication_mult_21_n43) );
  XOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U42 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_13__9_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_13__10_), .Z(
        my_filter_adder_mult_1_multiplication_mult_21_n42) );
  XOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U36 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_13__5_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_13__6_), .Z(
        my_filter_adder_mult_1_multiplication_mult_21_n36) );
  XOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U35 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_13__3_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_13__4_), .Z(
        my_filter_adder_mult_1_multiplication_mult_21_n35) );
  XOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U34 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_13__1_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_13__2_), .Z(
        my_filter_adder_mult_1_multiplication_mult_21_n34) );
  XOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U32 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_13__6_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_13__7_), .Z(
        my_filter_adder_mult_1_multiplication_mult_21_n32) );
  XOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U31 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_13__4_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_13__5_), .Z(
        my_filter_adder_mult_1_multiplication_mult_21_n31) );
  XOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U30 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_13__2_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_13__3_), .Z(
        my_filter_adder_mult_1_multiplication_mult_21_n30) );
  XOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U29 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_13__0_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_13__1_), .Z(
        my_filter_adder_mult_1_multiplication_mult_21_n29) );
  XOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U27 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_1__1_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_ab_0__2_), .Z(
        my_filter_adder_mult_1_multiplication_mult_21_n28) );
  XOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U26 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_13__12_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_13__13_), .Z(
        my_filter_adder_mult_1_multiplication_mult_21_n27) );
  XOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U25 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_1__12_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_ab_0__13_), .Z(
        my_filter_adder_mult_1_multiplication_mult_21_n26) );
  XOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U24 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_1__2_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_ab_0__3_), .Z(
        my_filter_adder_mult_1_multiplication_mult_21_n25) );
  XOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U23 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_1__3_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_ab_0__4_), .Z(
        my_filter_adder_mult_1_multiplication_mult_21_n24) );
  XOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U22 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_1__4_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_ab_0__5_), .Z(
        my_filter_adder_mult_1_multiplication_mult_21_n23) );
  XOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U21 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_1__5_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_ab_0__6_), .Z(
        my_filter_adder_mult_1_multiplication_mult_21_n22) );
  XOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U20 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_1__6_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_ab_0__7_), .Z(
        my_filter_adder_mult_1_multiplication_mult_21_n21) );
  XOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U19 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_1__7_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_ab_0__8_), .Z(
        my_filter_adder_mult_1_multiplication_mult_21_n20) );
  XOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U18 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_1__8_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_ab_0__9_), .Z(
        my_filter_adder_mult_1_multiplication_mult_21_n19) );
  XOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U17 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_1__9_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_ab_0__10_), .Z(
        my_filter_adder_mult_1_multiplication_mult_21_n18) );
  XOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U16 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_1__10_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_ab_0__11_), .Z(
        my_filter_adder_mult_1_multiplication_mult_21_n17) );
  XOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_U15 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_1__11_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_ab_0__12_), .Z(
        my_filter_adder_mult_1_multiplication_mult_21_n16) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S3_2_12 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_2__12_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_n15), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_ab_1__13_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_2__12_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_2__12_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_2_11 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_2__11_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_n4), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_n26), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_2__11_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_2__11_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_2_10 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_2__10_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_n5), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_n16), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_2__10_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_2__10_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_2_9 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_2__9_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_n6), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_n17), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_2__9_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_2__9_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_2_8 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_2__8_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_n7), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_n18), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_2__8_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_2__8_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_2_7 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_2__7_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_n8), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_n19), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_2__7_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_2__7_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_2_6 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_2__6_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_n9), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_n20), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_2__6_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_2__6_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_2_5 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_2__5_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_n10), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_n21), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_2__5_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_2__5_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_2_4 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_2__4_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_n11), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_n22), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_2__4_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_2__4_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_2_3 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_2__3_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_n12), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_n23), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_2__3_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_2__3_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_2_2 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_2__2_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_n13), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_n24), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_2__2_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_2__2_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_2_1 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_2__1_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_n14), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_n25), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_2__1_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_2__1_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S1_2_0 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_2__0_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_1__0_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_n28), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_2__0_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_A1_0_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S3_3_12 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_3__12_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_2__12_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_ab_2__13_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_3__12_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_3__12_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_3_11 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_3__11_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_2__11_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_2__12_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_3__11_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_3__11_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_3_10 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_3__10_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_2__10_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_2__11_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_3__10_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_3__10_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_3_9 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_3__9_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_2__9_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_2__10_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_3__9_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_3__9_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_3_8 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_3__8_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_2__8_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_2__9_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_3__8_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_3__8_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_3_7 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_3__7_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_2__7_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_2__8_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_3__7_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_3__7_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_3_6 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_3__6_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_2__6_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_2__7_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_3__6_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_3__6_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_3_5 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_3__5_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_2__5_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_2__6_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_3__5_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_3__5_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_3_4 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_3__4_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_2__4_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_2__5_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_3__4_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_3__4_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_3_3 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_3__3_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_2__3_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_2__4_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_3__3_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_3__3_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_3_2 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_3__2_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_2__2_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_2__3_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_3__2_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_3__2_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_3_1 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_3__1_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_2__1_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_2__2_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_3__1_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_3__1_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S1_3_0 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_3__0_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_2__0_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_2__1_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_3__0_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_A1_1_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S3_4_12 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_4__12_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_3__12_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_ab_3__13_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_4__12_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_4__12_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_4_11 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_4__11_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_3__11_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_3__12_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_4__11_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_4__11_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_4_10 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_4__10_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_3__10_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_3__11_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_4__10_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_4__10_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_4_9 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_4__9_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_3__9_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_3__10_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_4__9_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_4__9_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_4_8 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_4__8_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_3__8_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_3__9_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_4__8_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_4__8_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_4_7 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_4__7_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_3__7_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_3__8_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_4__7_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_4__7_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_4_6 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_4__6_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_3__6_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_3__7_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_4__6_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_4__6_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_4_5 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_4__5_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_3__5_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_3__6_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_4__5_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_4__5_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_4_4 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_4__4_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_3__4_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_3__5_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_4__4_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_4__4_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_4_3 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_4__3_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_3__3_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_3__4_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_4__3_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_4__3_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_4_2 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_4__2_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_3__2_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_3__3_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_4__2_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_4__2_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_4_1 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_4__1_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_3__1_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_3__2_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_4__1_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_4__1_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S1_4_0 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_4__0_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_3__0_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_3__1_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_4__0_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_A1_2_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S3_5_12 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_5__12_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_4__12_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_ab_4__13_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_5__12_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_5__12_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_5_11 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_5__11_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_4__11_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_4__12_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_5__11_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_5__11_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_5_10 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_5__10_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_4__10_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_4__11_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_5__10_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_5__10_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_5_9 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_5__9_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_4__9_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_4__10_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_5__9_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_5__9_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_5_8 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_5__8_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_4__8_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_4__9_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_5__8_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_5__8_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_5_7 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_5__7_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_4__7_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_4__8_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_5__7_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_5__7_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_5_6 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_5__6_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_4__6_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_4__7_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_5__6_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_5__6_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_5_5 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_5__5_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_4__5_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_4__6_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_5__5_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_5__5_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_5_4 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_5__4_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_4__4_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_4__5_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_5__4_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_5__4_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_5_3 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_5__3_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_4__3_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_4__4_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_5__3_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_5__3_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_5_2 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_5__2_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_4__2_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_4__3_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_5__2_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_5__2_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_5_1 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_5__1_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_4__1_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_4__2_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_5__1_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_5__1_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S1_5_0 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_5__0_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_4__0_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_4__1_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_5__0_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_A1_3_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S3_6_12 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_6__12_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_5__12_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_ab_5__13_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_6__12_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_6__12_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_6_11 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_6__11_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_5__11_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_5__12_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_6__11_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_6__11_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_6_10 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_6__10_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_5__10_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_5__11_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_6__10_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_6__10_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_6_9 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_6__9_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_5__9_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_5__10_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_6__9_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_6__9_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_6_8 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_6__8_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_5__8_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_5__9_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_6__8_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_6__8_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_6_7 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_6__7_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_5__7_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_5__8_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_6__7_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_6__7_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_6_6 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_6__6_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_5__6_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_5__7_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_6__6_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_6__6_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_6_5 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_6__5_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_5__5_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_5__6_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_6__5_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_6__5_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_6_4 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_6__4_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_5__4_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_5__5_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_6__4_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_6__4_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_6_3 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_6__3_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_5__3_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_5__4_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_6__3_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_6__3_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_6_2 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_6__2_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_5__2_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_5__3_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_6__2_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_6__2_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_6_1 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_6__1_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_5__1_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_5__2_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_6__1_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_6__1_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S1_6_0 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_6__0_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_5__0_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_5__1_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_6__0_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_A1_4_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S3_7_12 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_7__12_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_6__12_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_ab_6__13_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_7__12_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_7__12_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_7_11 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_7__11_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_6__11_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_6__12_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_7__11_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_7__11_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_7_10 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_7__10_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_6__10_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_6__11_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_7__10_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_7__10_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_7_9 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_7__9_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_6__9_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_6__10_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_7__9_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_7__9_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_7_8 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_7__8_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_6__8_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_6__9_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_7__8_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_7__8_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_7_7 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_7__7_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_6__7_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_6__8_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_7__7_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_7__7_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_7_6 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_7__6_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_6__6_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_6__7_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_7__6_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_7__6_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_7_5 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_7__5_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_6__5_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_6__6_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_7__5_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_7__5_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_7_4 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_7__4_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_6__4_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_6__5_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_7__4_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_7__4_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_7_3 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_7__3_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_6__3_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_6__4_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_7__3_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_7__3_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_7_2 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_7__2_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_6__2_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_6__3_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_7__2_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_7__2_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_7_1 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_7__1_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_6__1_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_6__2_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_7__1_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_7__1_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S1_7_0 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_7__0_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_6__0_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_6__1_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_7__0_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_A1_5_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S3_8_12 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_8__12_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_7__12_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_ab_7__13_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_8__12_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_8__12_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_8_11 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_8__11_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_7__11_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_7__12_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_8__11_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_8__11_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_8_10 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_8__10_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_7__10_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_7__11_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_8__10_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_8__10_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_8_9 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_8__9_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_7__9_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_7__10_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_8__9_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_8__9_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_8_8 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_8__8_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_7__8_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_7__9_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_8__8_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_8__8_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_8_7 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_8__7_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_7__7_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_7__8_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_8__7_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_8__7_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_8_6 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_8__6_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_7__6_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_7__7_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_8__6_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_8__6_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_8_5 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_8__5_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_7__5_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_7__6_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_8__5_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_8__5_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_8_4 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_8__4_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_7__4_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_7__5_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_8__4_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_8__4_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_8_3 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_8__3_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_7__3_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_7__4_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_8__3_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_8__3_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_8_2 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_8__2_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_7__2_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_7__3_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_8__2_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_8__2_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_8_1 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_8__1_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_7__1_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_7__2_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_8__1_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_8__1_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S1_8_0 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_8__0_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_7__0_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_7__1_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_8__0_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_A1_6_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S3_9_12 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_9__12_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_8__12_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_ab_8__13_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_9__12_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_9__12_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_9_11 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_9__11_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_8__11_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_8__12_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_9__11_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_9__11_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_9_10 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_9__10_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_8__10_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_8__11_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_9__10_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_9__10_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_9_9 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_9__9_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_8__9_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_8__10_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_9__9_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_9__9_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_9_8 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_9__8_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_8__8_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_8__9_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_9__8_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_9__8_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_9_7 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_9__7_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_8__7_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_8__8_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_9__7_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_9__7_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_9_6 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_9__6_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_8__6_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_8__7_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_9__6_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_9__6_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_9_5 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_9__5_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_8__5_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_8__6_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_9__5_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_9__5_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_9_4 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_9__4_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_8__4_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_8__5_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_9__4_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_9__4_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_9_3 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_9__3_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_8__3_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_8__4_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_9__3_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_9__3_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_9_2 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_9__2_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_8__2_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_8__3_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_9__2_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_9__2_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_9_1 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_9__1_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_8__1_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_8__2_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_9__1_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_9__1_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S1_9_0 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_9__0_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_8__0_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_8__1_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_9__0_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_A1_7_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S3_10_12 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_10__12_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_9__12_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_ab_9__13_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_10__12_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_10__12_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_10_11 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_10__11_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_9__11_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_9__12_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_10__11_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_10__11_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_10_10 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_10__10_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_9__10_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_9__11_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_10__10_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_10__10_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_10_9 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_10__9_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_9__9_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_9__10_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_10__9_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_10__9_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_10_8 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_10__8_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_9__8_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_9__9_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_10__8_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_10__8_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_10_7 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_10__7_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_9__7_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_9__8_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_10__7_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_10__7_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_10_6 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_10__6_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_9__6_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_9__7_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_10__6_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_10__6_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_10_5 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_10__5_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_9__5_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_9__6_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_10__5_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_10__5_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_10_4 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_10__4_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_9__4_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_9__5_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_10__4_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_10__4_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_10_3 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_10__3_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_9__3_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_9__4_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_10__3_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_10__3_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_10_2 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_10__2_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_9__2_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_9__3_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_10__2_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_10__2_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_10_1 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_10__1_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_9__1_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_9__2_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_10__1_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_10__1_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S1_10_0 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_10__0_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_9__0_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_9__1_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_10__0_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_A1_8_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S3_11_12 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_11__12_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_10__12_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_ab_10__13_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_11__12_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_11__12_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_11_11 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_11__11_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_10__11_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_10__12_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_11__11_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_11__11_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_11_10 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_11__10_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_10__10_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_10__11_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_11__10_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_11__10_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_11_9 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_11__9_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_10__9_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_10__10_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_11__9_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_11__9_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_11_8 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_11__8_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_10__8_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_10__9_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_11__8_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_11__8_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_11_7 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_11__7_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_10__7_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_10__8_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_11__7_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_11__7_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_11_6 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_11__6_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_10__6_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_10__7_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_11__6_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_11__6_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_11_5 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_11__5_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_10__5_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_10__6_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_11__5_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_11__5_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_11_4 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_11__4_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_10__4_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_10__5_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_11__4_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_11__4_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_11_3 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_11__3_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_10__3_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_10__4_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_11__3_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_11__3_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_11_2 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_11__2_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_10__2_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_10__3_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_11__2_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_11__2_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_11_1 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_11__1_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_10__1_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_10__2_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_11__1_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_11__1_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S1_11_0 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_11__0_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_10__0_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_10__1_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_11__0_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_A1_9_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S3_12_12 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_12__12_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_11__12_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_ab_11__13_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_12__12_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_12__12_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_12_11 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_12__11_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_11__11_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_11__12_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_12__11_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_12__11_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_12_10 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_12__10_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_11__10_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_11__11_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_12__10_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_12__10_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_12_9 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_12__9_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_11__9_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_11__10_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_12__9_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_12__9_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_12_8 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_12__8_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_11__8_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_11__9_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_12__8_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_12__8_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_12_7 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_12__7_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_11__7_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_11__8_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_12__7_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_12__7_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_12_6 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_12__6_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_11__6_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_11__7_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_12__6_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_12__6_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_12_5 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_12__5_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_11__5_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_11__6_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_12__5_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_12__5_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_12_4 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_12__4_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_11__4_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_11__5_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_12__4_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_12__4_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_12_3 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_12__3_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_11__3_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_11__4_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_12__3_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_12__3_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_12_2 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_12__2_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_11__2_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_11__3_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_12__2_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_12__2_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S2_12_1 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_12__1_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_11__1_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_11__2_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_12__1_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_12__1_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S1_12_0 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_12__0_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_11__0_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_11__1_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_12__0_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_A1_10_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S14_13 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_n86), .B(
        my_filter_adder_mult_1_multiplication_mult_21_n100), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_ab_13__13_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_13__13_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_13__13_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S5_12 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_13__12_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_12__12_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_ab_12__13_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_13__12_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_13__12_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S4_11 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_13__11_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_12__11_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_12__12_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_13__11_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_13__11_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S4_10 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_13__10_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_12__10_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_12__11_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_13__10_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_13__10_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S4_9 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_13__9_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_12__9_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_12__10_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_13__9_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_13__9_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S4_8 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_13__8_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_12__8_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_12__9_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_13__8_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_13__8_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S4_7 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_13__7_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_12__7_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_12__8_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_13__7_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_13__7_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S4_6 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_13__6_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_12__6_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_12__7_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_13__6_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_13__6_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S4_5 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_13__5_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_12__5_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_12__6_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_13__5_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_13__5_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S4_4 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_13__4_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_12__4_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_12__5_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_13__4_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_13__4_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S4_3 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_13__3_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_12__3_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_12__4_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_13__3_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_13__3_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S4_2 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_13__2_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_12__2_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_12__3_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_13__2_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_13__2_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S4_1 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_13__1_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_12__1_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_12__2_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_13__1_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_13__1_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S4_0 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_ab_13__0_), .B(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_12__0_), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_12__1_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_CARRYB_13__0_), .S(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_13__0_) );
  FA_X1 my_filter_adder_mult_1_multiplication_mult_21_S14_13_0 ( .A(
        my_filter_q_reg_chain_2__13_), .B(my_filter_q_reg_coeff[125]), .CI(
        my_filter_adder_mult_1_multiplication_mult_21_SUMB_13__0_), .CO(
        my_filter_adder_mult_1_multiplication_mult_21_A2_12_), .S(
        my_filter_adder_mult_1_res_mult[0]) );
  NAND2_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U72 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_A2_12_), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n29), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n56) );
  OAI21_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U71 ( .B1(
        my_filter_adder_mult_1_multiplication_mult_21_A2_12_), .B2(
        my_filter_adder_mult_1_multiplication_mult_21_n29), .A(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n56), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n59) );
  INV_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U70 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n59), .ZN(
        my_filter_adder_mult_1_res_mult[1]) );
  OAI21_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U69 ( .B1(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n15), .B2(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n16), .A(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n17), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n13) );
  AND2_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U68 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n51), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n49), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n20) );
  AND2_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U66 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n50), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n43), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n28) );
  AND2_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U65 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n41), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n32), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n36) );
  NAND2_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U64 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n47), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n44), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n17) );
  NAND2_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U63 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n46), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n42), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n25) );
  NAND2_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U61 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n45), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n48), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n33) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U60 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n47), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n44), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n15) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U59 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n46), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n42), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n23) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U58 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n45), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n48), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n31) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U56 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n51), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n49), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n21) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U55 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n50), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n43), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n29) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U54 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n41), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n32), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n37) );
  AND2_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U53 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n33), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n31), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n44) );
  AND2_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U51 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n40), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n30), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n52) );
  NAND2_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U50 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n39), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n36), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n41) );
  NAND2_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U49 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n38), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n35), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n49) );
  NAND2_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U48 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n37), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n34), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n57) );
  INV_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U46 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n55), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n60) );
  NAND2_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U45 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n60), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n57), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n58) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U44 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n39), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n36), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n39) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U43 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n38), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n35), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n47) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U41 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n37), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n34), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n55) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U40 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n33), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n31), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n45) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U39 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_n40), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_n30), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n53) );
  OAI21_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U38 ( .B1(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n55), .B2(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n56), .A(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n57), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n51) );
  INV_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U36 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n15), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n62) );
  NAND2_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U35 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n62), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n17), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n18) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U34 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n20), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n21), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n22) );
  INV_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U33 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n23), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n64) );
  NAND2_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U31 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n64), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n25), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n26) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U30 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n28), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n29), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n30) );
  INV_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U29 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n31), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n70) );
  NAND2_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U28 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n70), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n33), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n34) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U26 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n36), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n37), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n38) );
  INV_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U25 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n39), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n68) );
  NAND2_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U24 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n68), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n41), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n42) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U23 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n44), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n45), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n46) );
  INV_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U21 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n47), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n66) );
  NAND2_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U20 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n66), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n49), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n50) );
  NOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U19 ( .A1(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n52), .A2(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n53), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n54) );
  OAI21_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U18 ( .B1(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n23), .B2(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n24), .A(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n25), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n19) );
  OAI21_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U16 ( .B1(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n31), .B2(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n32), .A(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n33), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n27) );
  OAI21_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U13 ( .B1(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n39), .B2(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n40), .A(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n41), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n35) );
  OAI21_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U12 ( .B1(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n47), .B2(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n48), .A(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n49), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n43) );
  INV_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U11 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n21), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n63) );
  AOI21_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U10 ( .B1(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n63), .B2(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n19), .A(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n20), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n16) );
  INV_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U9 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n29), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n71) );
  AOI21_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U8 ( .B1(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n71), .B2(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n27), .A(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n28), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n24) );
  INV_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U7 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n37), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n69) );
  AOI21_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U6 ( .B1(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n69), .B2(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n35), .A(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n36), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n32) );
  INV_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U5 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n45), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n67) );
  AOI21_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U4 ( .B1(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n67), .B2(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n43), .A(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n44), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n40) );
  INV_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U3 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n53), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n65) );
  AOI21_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U2 ( .B1(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n65), .B2(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n51), .A(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n52), .ZN(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n48) );
  XOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U67 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n56), .B(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n58), .Z(
        my_filter_adder_mult_1_res_mult[2]) );
  XOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U62 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n51), .B(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n54), .Z(
        my_filter_adder_mult_1_res_mult[3]) );
  XOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U57 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n50), .B(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n48), .Z(
        my_filter_adder_mult_1_res_mult[4]) );
  XOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U52 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n43), .B(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n46), .Z(
        my_filter_adder_mult_1_res_mult[5]) );
  XOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U47 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n42), .B(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n40), .Z(
        my_filter_adder_mult_1_res_mult[6]) );
  XOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U42 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n35), .B(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n38), .Z(
        my_filter_adder_mult_1_res_mult[7]) );
  XOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U37 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n34), .B(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n32), .Z(
        my_filter_adder_mult_1_res_mult[8]) );
  XOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U32 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n27), .B(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n30), .Z(
        my_filter_adder_mult_1_res_mult[9]) );
  XOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U27 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n26), .B(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n24), .Z(
        my_filter_adder_mult_1_res_mult[10]) );
  XOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U22 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n19), .B(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n22), .Z(
        my_filter_adder_mult_1_res_mult[11]) );
  XOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U17 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n18), .B(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n16), .Z(
        my_filter_adder_mult_1_res_mult[12]) );
  XOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U15 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_n52), .B(
        my_filter_adder_mult_1_multiplication_mult_21_n27), .Z(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n14) );
  XOR2_X1 my_filter_adder_mult_1_multiplication_mult_21_FS_1_U14 ( .A(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n13), .B(
        my_filter_adder_mult_1_multiplication_mult_21_FS_1_n14), .Z(
        my_filter_adder_mult_1_res_mult[13]) );
  AND2_X1 my_filter_adder_mult_1_addition_add_19_U1 ( .A1(
        my_filter_data_sum[126]), .A2(my_filter_adder_mult_1_res_mult[0]), 
        .ZN(my_filter_adder_mult_1_addition_add_19_n1) );
  XOR2_X1 my_filter_adder_mult_1_addition_add_19_U2 ( .A(
        my_filter_data_sum[126]), .B(my_filter_adder_mult_1_res_mult[0]), .Z(
        my_filter_data_sum[112]) );
  FA_X1 my_filter_adder_mult_1_addition_add_19_U1_1 ( .A(
        my_filter_adder_mult_1_res_mult[1]), .B(my_filter_data_sum[127]), .CI(
        my_filter_adder_mult_1_addition_add_19_n1), .CO(
        my_filter_adder_mult_1_addition_add_19_carry[2]), .S(
        my_filter_data_sum[113]) );
  FA_X1 my_filter_adder_mult_1_addition_add_19_U1_2 ( .A(
        my_filter_adder_mult_1_res_mult[2]), .B(my_filter_data_sum[128]), .CI(
        my_filter_adder_mult_1_addition_add_19_carry[2]), .CO(
        my_filter_adder_mult_1_addition_add_19_carry[3]), .S(
        my_filter_data_sum[114]) );
  FA_X1 my_filter_adder_mult_1_addition_add_19_U1_3 ( .A(
        my_filter_adder_mult_1_res_mult[3]), .B(my_filter_data_sum[129]), .CI(
        my_filter_adder_mult_1_addition_add_19_carry[3]), .CO(
        my_filter_adder_mult_1_addition_add_19_carry[4]), .S(
        my_filter_data_sum[115]) );
  FA_X1 my_filter_adder_mult_1_addition_add_19_U1_4 ( .A(
        my_filter_adder_mult_1_res_mult[4]), .B(my_filter_data_sum[130]), .CI(
        my_filter_adder_mult_1_addition_add_19_carry[4]), .CO(
        my_filter_adder_mult_1_addition_add_19_carry[5]), .S(
        my_filter_data_sum[116]) );
  FA_X1 my_filter_adder_mult_1_addition_add_19_U1_5 ( .A(
        my_filter_adder_mult_1_res_mult[5]), .B(my_filter_data_sum[131]), .CI(
        my_filter_adder_mult_1_addition_add_19_carry[5]), .CO(
        my_filter_adder_mult_1_addition_add_19_carry[6]), .S(
        my_filter_data_sum[117]) );
  FA_X1 my_filter_adder_mult_1_addition_add_19_U1_6 ( .A(
        my_filter_adder_mult_1_res_mult[6]), .B(my_filter_data_sum[132]), .CI(
        my_filter_adder_mult_1_addition_add_19_carry[6]), .CO(
        my_filter_adder_mult_1_addition_add_19_carry[7]), .S(
        my_filter_data_sum[118]) );
  FA_X1 my_filter_adder_mult_1_addition_add_19_U1_7 ( .A(
        my_filter_adder_mult_1_res_mult[7]), .B(my_filter_data_sum[133]), .CI(
        my_filter_adder_mult_1_addition_add_19_carry[7]), .CO(
        my_filter_adder_mult_1_addition_add_19_carry[8]), .S(
        my_filter_data_sum[119]) );
  FA_X1 my_filter_adder_mult_1_addition_add_19_U1_8 ( .A(
        my_filter_adder_mult_1_res_mult[8]), .B(my_filter_data_sum[134]), .CI(
        my_filter_adder_mult_1_addition_add_19_carry[8]), .CO(
        my_filter_adder_mult_1_addition_add_19_carry[9]), .S(
        my_filter_data_sum[120]) );
  FA_X1 my_filter_adder_mult_1_addition_add_19_U1_9 ( .A(
        my_filter_adder_mult_1_res_mult[9]), .B(my_filter_data_sum[135]), .CI(
        my_filter_adder_mult_1_addition_add_19_carry[9]), .CO(
        my_filter_adder_mult_1_addition_add_19_carry[10]), .S(
        my_filter_data_sum[121]) );
  FA_X1 my_filter_adder_mult_1_addition_add_19_U1_10 ( .A(
        my_filter_adder_mult_1_res_mult[10]), .B(my_filter_data_sum[136]), 
        .CI(my_filter_adder_mult_1_addition_add_19_carry[10]), .CO(
        my_filter_adder_mult_1_addition_add_19_carry[11]), .S(
        my_filter_data_sum[122]) );
  FA_X1 my_filter_adder_mult_1_addition_add_19_U1_11 ( .A(
        my_filter_adder_mult_1_res_mult[11]), .B(my_filter_data_sum[137]), 
        .CI(my_filter_adder_mult_1_addition_add_19_carry[11]), .CO(
        my_filter_adder_mult_1_addition_add_19_carry[12]), .S(
        my_filter_data_sum[123]) );
  FA_X1 my_filter_adder_mult_1_addition_add_19_U1_12 ( .A(
        my_filter_adder_mult_1_res_mult[12]), .B(my_filter_data_sum[138]), 
        .CI(my_filter_adder_mult_1_addition_add_19_carry[12]), .CO(
        my_filter_adder_mult_1_addition_add_19_carry[13]), .S(
        my_filter_data_sum[124]) );
  FA_X1 my_filter_adder_mult_1_addition_add_19_U1_13 ( .A(
        my_filter_adder_mult_1_res_mult[13]), .B(my_filter_data_sum[139]), 
        .CI(my_filter_adder_mult_1_addition_add_19_carry[13]), .S(
        my_filter_data_sum[125]) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U276 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_12__12_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U275 ( .A1(
        my_filter_q_reg_chain_3__11_), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_11__13_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U274 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_11__12_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U273 ( .A1(
        my_filter_q_reg_chain_3__10_), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_10__13_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U272 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_10__12_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U271 ( .A1(
        my_filter_q_reg_chain_3__9_), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_9__13_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U270 ( .A1(
        my_filter_q_reg_chain_3__8_), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_8__13_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U269 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n101), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_9__12_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U268 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_8__12_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U267 ( .A1(
        my_filter_q_reg_chain_3__7_), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_7__13_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U266 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_7__12_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U265 ( .A1(
        my_filter_q_reg_chain_3__6_), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_6__13_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U264 ( .A1(
        my_filter_q_reg_coeff[108]), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_13__10_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U263 ( .A1(
        my_filter_q_reg_coeff[109]), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_13__11_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U262 ( .A1(
        my_filter_q_reg_coeff[106]), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_13__8_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U261 ( .A1(
        my_filter_q_reg_coeff[107]), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_13__9_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U260 ( .A1(
        my_filter_q_reg_coeff[104]), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_13__6_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U259 ( .A1(
        my_filter_q_reg_coeff[105]), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_13__7_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U258 ( .A1(
        my_filter_q_reg_coeff[110]), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_13__12_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U257 ( .A1(
        my_filter_q_reg_chain_3__12_), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_12__13_) );
  INV_X1 my_filter_adder_mult_2_multiplication_mult_21_U256 ( .A(
        my_filter_q_reg_chain_3__9_), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_n90) );
  INV_X1 my_filter_adder_mult_2_multiplication_mult_21_U255 ( .A(
        my_filter_q_reg_chain_3__12_), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_n87) );
  INV_X1 my_filter_adder_mult_2_multiplication_mult_21_U254 ( .A(
        my_filter_q_reg_chain_3__11_), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_n88) );
  INV_X1 my_filter_adder_mult_2_multiplication_mult_21_U253 ( .A(
        my_filter_q_reg_chain_3__10_), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_n89) );
  INV_X1 my_filter_adder_mult_2_multiplication_mult_21_U252 ( .A(
        my_filter_q_reg_chain_3__8_), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_n91) );
  INV_X1 my_filter_adder_mult_2_multiplication_mult_21_U251 ( .A(
        my_filter_q_reg_chain_3__7_), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_n92) );
  INV_X1 my_filter_adder_mult_2_multiplication_mult_21_U250 ( .A(
        my_filter_q_reg_chain_3__6_), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_n93) );
  INV_X1 my_filter_adder_mult_2_multiplication_mult_21_U249 ( .A(
        my_filter_q_reg_chain_3__13_), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_n86) );
  AND2_X1 my_filter_adder_mult_2_multiplication_mult_21_U248 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_ab_0__13_), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_ab_1__12_), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_n15) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U247 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_2__12_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U246 ( .A1(
        my_filter_q_reg_chain_3__1_), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_1__13_) );
  AND3_X1 my_filter_adder_mult_2_multiplication_mult_21_U245 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_ab_1__1_), .A2(
        my_filter_q_reg_coeff[98]), .A3(my_filter_q_reg_chain_3__0_), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_1__0_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U244 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_12__0_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U243 ( .A1(
        my_filter_q_reg_coeff[98]), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_13__0_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U242 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_6__12_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U241 ( .A1(
        my_filter_q_reg_chain_3__5_), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_5__13_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U240 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_5__12_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U239 ( .A1(
        my_filter_q_reg_chain_3__4_), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_4__13_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U238 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_4__12_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U237 ( .A1(
        my_filter_q_reg_chain_3__3_), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_3__13_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U236 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_3__12_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U235 ( .A1(
        my_filter_q_reg_chain_3__2_), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_2__13_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U234 ( .A1(
        my_filter_q_reg_coeff[102]), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_13__4_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U233 ( .A1(
        my_filter_q_reg_coeff[103]), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_13__5_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U232 ( .A1(
        my_filter_q_reg_coeff[99]), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_13__1_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U231 ( .A1(
        my_filter_q_reg_coeff[100]), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_13__2_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U230 ( .A1(
        my_filter_q_reg_coeff[101]), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_13__3_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U229 ( .A1(
        my_filter_q_reg_chain_3__0_), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_0__13_) );
  INV_X1 my_filter_adder_mult_2_multiplication_mult_21_U228 ( .A(
        my_filter_q_reg_coeff[111]), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_n100) );
  INV_X1 my_filter_adder_mult_2_multiplication_mult_21_U227 ( .A(
        my_filter_q_reg_coeff[98]), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_n113) );
  INV_X1 my_filter_adder_mult_2_multiplication_mult_21_U226 ( .A(
        my_filter_q_reg_chain_3__0_), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_n99) );
  INV_X1 my_filter_adder_mult_2_multiplication_mult_21_U225 ( .A(
        my_filter_q_reg_coeff[99]), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_n112) );
  INV_X1 my_filter_adder_mult_2_multiplication_mult_21_U224 ( .A(
        my_filter_q_reg_chain_3__1_), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_n98) );
  INV_X1 my_filter_adder_mult_2_multiplication_mult_21_U223 ( .A(
        my_filter_q_reg_coeff[110]), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_n101) );
  INV_X1 my_filter_adder_mult_2_multiplication_mult_21_U222 ( .A(
        my_filter_q_reg_coeff[108]), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_n103) );
  INV_X1 my_filter_adder_mult_2_multiplication_mult_21_U221 ( .A(
        my_filter_q_reg_coeff[109]), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_n102) );
  INV_X1 my_filter_adder_mult_2_multiplication_mult_21_U220 ( .A(
        my_filter_q_reg_coeff[106]), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_n105) );
  INV_X1 my_filter_adder_mult_2_multiplication_mult_21_U219 ( .A(
        my_filter_q_reg_coeff[107]), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_n104) );
  INV_X1 my_filter_adder_mult_2_multiplication_mult_21_U218 ( .A(
        my_filter_q_reg_coeff[103]), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_n108) );
  INV_X1 my_filter_adder_mult_2_multiplication_mult_21_U217 ( .A(
        my_filter_q_reg_coeff[104]), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_n107) );
  INV_X1 my_filter_adder_mult_2_multiplication_mult_21_U216 ( .A(
        my_filter_q_reg_coeff[105]), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_n106) );
  INV_X1 my_filter_adder_mult_2_multiplication_mult_21_U215 ( .A(
        my_filter_q_reg_coeff[100]), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_n111) );
  INV_X1 my_filter_adder_mult_2_multiplication_mult_21_U214 ( .A(
        my_filter_q_reg_coeff[101]), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_n110) );
  INV_X1 my_filter_adder_mult_2_multiplication_mult_21_U213 ( .A(
        my_filter_q_reg_coeff[102]), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_n109) );
  INV_X1 my_filter_adder_mult_2_multiplication_mult_21_U212 ( .A(
        my_filter_q_reg_chain_3__5_), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_n94) );
  INV_X1 my_filter_adder_mult_2_multiplication_mult_21_U211 ( .A(
        my_filter_q_reg_chain_3__4_), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_n95) );
  INV_X1 my_filter_adder_mult_2_multiplication_mult_21_U210 ( .A(
        my_filter_q_reg_chain_3__2_), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_n97) );
  INV_X1 my_filter_adder_mult_2_multiplication_mult_21_U209 ( .A(
        my_filter_q_reg_chain_3__3_), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_n96) );
  AND2_X1 my_filter_adder_mult_2_multiplication_mult_21_U208 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_13__12_), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_13__13_), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_n3) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U207 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n100), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_13__13_) );
  AND2_X1 my_filter_adder_mult_2_multiplication_mult_21_U206 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_13__11_), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_13__12_), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_n52) );
  AND2_X1 my_filter_adder_mult_2_multiplication_mult_21_U205 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_13__9_), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_13__10_), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_n50) );
  AND2_X1 my_filter_adder_mult_2_multiplication_mult_21_U204 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_13__7_), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_13__8_), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_n49) );
  AND2_X1 my_filter_adder_mult_2_multiplication_mult_21_U203 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_13__5_), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_13__6_), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_n48) );
  AND2_X1 my_filter_adder_mult_2_multiplication_mult_21_U202 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_13__10_), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_13__11_), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_n45) );
  AND2_X1 my_filter_adder_mult_2_multiplication_mult_21_U201 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_13__8_), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_13__9_), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_n44) );
  AND2_X1 my_filter_adder_mult_2_multiplication_mult_21_U200 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_13__6_), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_13__7_), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_n43) );
  AND2_X1 my_filter_adder_mult_2_multiplication_mult_21_U199 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_13__4_), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_13__5_), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_n46) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U198 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_12__11_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U197 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_12__9_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U196 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_12__10_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U195 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_11__10_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U194 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_11__11_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U193 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_12__7_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U192 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_12__8_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U191 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_10__11_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U190 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_11__8_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U189 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_11__9_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U188 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_10__9_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U187 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_10__10_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U186 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n103), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_9__10_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U185 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n102), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_9__11_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U184 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_8__11_) );
  AND2_X1 my_filter_adder_mult_2_multiplication_mult_21_U183 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_13__3_), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_13__4_), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_n31) );
  AND2_X1 my_filter_adder_mult_2_multiplication_mult_21_U182 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_13__1_), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_13__2_), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_n37) );
  AND2_X1 my_filter_adder_mult_2_multiplication_mult_21_U181 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_13__2_), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_13__3_), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_n36) );
  AND2_X1 my_filter_adder_mult_2_multiplication_mult_21_U180 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_13__0_), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_13__1_), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_n35) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U179 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_12__1_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U178 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_10__0_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U177 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_11__0_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U176 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_11__1_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U175 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_10__1_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U174 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_8__0_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U173 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n113), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_9__0_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U172 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n112), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_9__1_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U171 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n110), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_9__3_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U170 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_8__1_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U169 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_8__3_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U168 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_6__0_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U167 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_7__0_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U166 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_7__1_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U165 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_7__3_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U164 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_7__4_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U163 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_7__5_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U162 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_6__1_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U161 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_6__3_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U160 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_6__5_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U159 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_4__0_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U158 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_5__0_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U157 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_5__1_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U156 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_5__3_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U155 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_5__4_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U154 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_5__5_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U153 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_5__6_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U152 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_5__7_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U151 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_4__1_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U150 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_4__3_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U149 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_4__5_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U148 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_2__0_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U147 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_3__0_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U146 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_3__1_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U145 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_3__3_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U144 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_3__4_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U143 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_3__5_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U142 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_3__6_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U141 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_3__7_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U140 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_3__8_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U139 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_3__9_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U138 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_12__5_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U137 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_12__6_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U136 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_11__6_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U135 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_11__7_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U134 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_12__2_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U133 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_12__3_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U132 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_12__4_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U131 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_10__7_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U130 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_10__8_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U129 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_11__3_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U128 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_11__4_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U127 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_11__5_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U126 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n105), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_9__8_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U125 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n104), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_9__9_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U124 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_10__4_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U123 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_10__5_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U122 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_10__6_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U121 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_8__9_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U120 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_8__10_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U119 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_11__2_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U118 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n108), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_9__5_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U117 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n107), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_9__6_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U116 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n106), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_9__7_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U115 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_7__10_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U114 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_7__11_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U113 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_10__2_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U112 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_10__3_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U111 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_8__6_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U110 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_8__7_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U109 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_8__8_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U108 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_6__11_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U107 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n111), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_9__2_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U106 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n109), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_9__4_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U105 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_7__7_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U104 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_7__8_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U103 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_7__9_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U102 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_8__2_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U101 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_8__4_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U100 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_8__5_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U99 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_6__8_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U98 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_6__9_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U97 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_6__10_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U96 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_7__2_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U95 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_7__6_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U94 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_5__9_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U93 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_5__10_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U92 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_5__11_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U91 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_6__2_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U90 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_6__4_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U89 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_6__6_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U88 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_6__7_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U87 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_4__10_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U86 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_4__11_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U85 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_5__2_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U84 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_5__8_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U83 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_3__11_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U82 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_4__2_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U81 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_4__4_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U80 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_4__6_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U79 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_4__7_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U78 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_4__8_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U77 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_4__9_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U76 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_3__2_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U75 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_3__10_) );
  AND2_X1 my_filter_adder_mult_2_multiplication_mult_21_U74 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_ab_0__2_), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_ab_1__1_), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_n14) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U73 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_2__1_) );
  AND2_X1 my_filter_adder_mult_2_multiplication_mult_21_U72 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_ab_0__3_), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_ab_1__2_), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_n13) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U71 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_2__2_) );
  AND2_X1 my_filter_adder_mult_2_multiplication_mult_21_U70 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_ab_0__4_), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_ab_1__3_), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_n12) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U69 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_2__3_) );
  AND2_X1 my_filter_adder_mult_2_multiplication_mult_21_U68 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_ab_0__5_), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_ab_1__4_), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_n11) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U67 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_2__4_) );
  AND2_X1 my_filter_adder_mult_2_multiplication_mult_21_U66 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_ab_0__6_), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_ab_1__5_), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_n10) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U65 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_2__5_) );
  AND2_X1 my_filter_adder_mult_2_multiplication_mult_21_U64 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_ab_0__7_), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_ab_1__6_), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_n9) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U63 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_2__6_) );
  AND2_X1 my_filter_adder_mult_2_multiplication_mult_21_U62 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_ab_0__8_), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_ab_1__7_), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_n8) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U61 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_2__7_) );
  AND2_X1 my_filter_adder_mult_2_multiplication_mult_21_U60 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_ab_0__9_), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_ab_1__8_), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_n7) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U59 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_2__8_) );
  AND2_X1 my_filter_adder_mult_2_multiplication_mult_21_U58 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_ab_0__10_), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_ab_1__9_), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_n6) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U57 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_2__9_) );
  AND2_X1 my_filter_adder_mult_2_multiplication_mult_21_U56 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_ab_0__11_), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_ab_1__10_), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_n5) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U55 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_2__10_) );
  AND2_X1 my_filter_adder_mult_2_multiplication_mult_21_U54 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_ab_0__12_), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_ab_1__11_), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_n4) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U52 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_2__11_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U50 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_1__12_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U49 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_1__2_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U48 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_1__3_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U46 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_1__4_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U45 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_1__5_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U44 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_1__6_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U43 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_1__7_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U37 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_1__8_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U36 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_1__9_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U35 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_1__10_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U31 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_1__11_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U14 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_0__2_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U13 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_0__3_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U12 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_0__4_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U11 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_0__5_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U10 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_0__6_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U9 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_0__7_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U8 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_0__8_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U7 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_0__9_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U6 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_0__10_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U5 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_0__11_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U4 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_0__12_) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U3 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n98), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n112), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_ab_1__1_) );
  INV_X1 my_filter_adder_mult_2_multiplication_mult_21_U2 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_13__13_), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_n85) );
  XOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U51 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_13__12_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_13__13_), .Z(
        my_filter_adder_mult_2_multiplication_mult_21_n51) );
  XOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U47 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_13__10_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_13__11_), .Z(
        my_filter_adder_mult_2_multiplication_mult_21_n47) );
  XOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U42 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_13__11_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_13__12_), .Z(
        my_filter_adder_mult_2_multiplication_mult_21_n42) );
  XOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U41 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_13__8_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_13__9_), .Z(
        my_filter_adder_mult_2_multiplication_mult_21_n41) );
  XOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U40 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_13__9_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_13__10_), .Z(
        my_filter_adder_mult_2_multiplication_mult_21_n40) );
  XOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U39 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_13__6_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_13__7_), .Z(
        my_filter_adder_mult_2_multiplication_mult_21_n39) );
  XOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U38 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_13__7_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_13__8_), .Z(
        my_filter_adder_mult_2_multiplication_mult_21_n38) );
  XOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U34 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_13__5_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_13__6_), .Z(
        my_filter_adder_mult_2_multiplication_mult_21_n34) );
  XOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U33 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_13__3_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_13__4_), .Z(
        my_filter_adder_mult_2_multiplication_mult_21_n33) );
  XOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U32 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_13__1_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_13__2_), .Z(
        my_filter_adder_mult_2_multiplication_mult_21_n32) );
  XOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U30 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_13__4_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_13__5_), .Z(
        my_filter_adder_mult_2_multiplication_mult_21_n30) );
  XOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U29 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_13__2_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_13__3_), .Z(
        my_filter_adder_mult_2_multiplication_mult_21_n29) );
  XOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U28 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_13__0_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_13__1_), .Z(
        my_filter_adder_mult_2_multiplication_mult_21_n28) );
  XOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U26 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_1__1_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_ab_0__2_), .Z(
        my_filter_adder_mult_2_multiplication_mult_21_n27) );
  XOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U25 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_1__12_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_ab_0__13_), .Z(
        my_filter_adder_mult_2_multiplication_mult_21_n26) );
  XOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U24 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_1__2_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_ab_0__3_), .Z(
        my_filter_adder_mult_2_multiplication_mult_21_n25) );
  XOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U23 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_1__3_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_ab_0__4_), .Z(
        my_filter_adder_mult_2_multiplication_mult_21_n24) );
  XOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U22 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_1__4_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_ab_0__5_), .Z(
        my_filter_adder_mult_2_multiplication_mult_21_n23) );
  XOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U21 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_1__5_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_ab_0__6_), .Z(
        my_filter_adder_mult_2_multiplication_mult_21_n22) );
  XOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U20 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_1__6_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_ab_0__7_), .Z(
        my_filter_adder_mult_2_multiplication_mult_21_n21) );
  XOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U19 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_1__7_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_ab_0__8_), .Z(
        my_filter_adder_mult_2_multiplication_mult_21_n20) );
  XOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U18 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_1__8_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_ab_0__9_), .Z(
        my_filter_adder_mult_2_multiplication_mult_21_n19) );
  XOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U17 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_1__9_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_ab_0__10_), .Z(
        my_filter_adder_mult_2_multiplication_mult_21_n18) );
  XOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U16 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_1__10_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_ab_0__11_), .Z(
        my_filter_adder_mult_2_multiplication_mult_21_n17) );
  XOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_U15 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_1__11_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_ab_0__12_), .Z(
        my_filter_adder_mult_2_multiplication_mult_21_n16) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S3_2_12 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_2__12_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_n15), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_ab_1__13_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_2__12_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_2__12_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_2_11 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_2__11_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_n4), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_n26), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_2__11_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_2__11_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_2_10 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_2__10_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_n5), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_n16), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_2__10_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_2__10_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_2_9 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_2__9_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_n6), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_n17), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_2__9_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_2__9_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_2_8 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_2__8_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_n7), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_n18), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_2__8_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_2__8_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_2_7 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_2__7_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_n8), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_n19), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_2__7_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_2__7_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_2_6 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_2__6_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_n9), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_n20), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_2__6_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_2__6_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_2_5 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_2__5_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_n10), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_n21), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_2__5_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_2__5_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_2_4 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_2__4_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_n11), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_n22), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_2__4_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_2__4_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_2_3 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_2__3_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_n12), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_n23), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_2__3_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_2__3_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_2_2 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_2__2_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_n13), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_n24), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_2__2_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_2__2_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_2_1 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_2__1_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_n14), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_n25), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_2__1_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_2__1_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S1_2_0 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_2__0_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_1__0_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_n27), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_2__0_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_A1_0_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S3_3_12 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_3__12_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_2__12_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_ab_2__13_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_3__12_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_3__12_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_3_11 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_3__11_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_2__11_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_2__12_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_3__11_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_3__11_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_3_10 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_3__10_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_2__10_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_2__11_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_3__10_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_3__10_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_3_9 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_3__9_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_2__9_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_2__10_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_3__9_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_3__9_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_3_8 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_3__8_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_2__8_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_2__9_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_3__8_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_3__8_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_3_7 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_3__7_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_2__7_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_2__8_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_3__7_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_3__7_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_3_6 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_3__6_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_2__6_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_2__7_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_3__6_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_3__6_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_3_5 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_3__5_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_2__5_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_2__6_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_3__5_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_3__5_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_3_4 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_3__4_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_2__4_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_2__5_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_3__4_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_3__4_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_3_3 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_3__3_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_2__3_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_2__4_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_3__3_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_3__3_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_3_2 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_3__2_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_2__2_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_2__3_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_3__2_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_3__2_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_3_1 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_3__1_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_2__1_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_2__2_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_3__1_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_3__1_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S1_3_0 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_3__0_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_2__0_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_2__1_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_3__0_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_A1_1_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S3_4_12 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_4__12_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_3__12_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_ab_3__13_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_4__12_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_4__12_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_4_11 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_4__11_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_3__11_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_3__12_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_4__11_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_4__11_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_4_10 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_4__10_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_3__10_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_3__11_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_4__10_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_4__10_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_4_9 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_4__9_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_3__9_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_3__10_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_4__9_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_4__9_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_4_8 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_4__8_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_3__8_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_3__9_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_4__8_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_4__8_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_4_7 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_4__7_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_3__7_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_3__8_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_4__7_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_4__7_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_4_6 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_4__6_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_3__6_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_3__7_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_4__6_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_4__6_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_4_5 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_4__5_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_3__5_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_3__6_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_4__5_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_4__5_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_4_4 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_4__4_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_3__4_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_3__5_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_4__4_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_4__4_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_4_3 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_4__3_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_3__3_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_3__4_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_4__3_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_4__3_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_4_2 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_4__2_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_3__2_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_3__3_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_4__2_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_4__2_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_4_1 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_4__1_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_3__1_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_3__2_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_4__1_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_4__1_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S1_4_0 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_4__0_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_3__0_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_3__1_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_4__0_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_A1_2_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S3_5_12 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_5__12_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_4__12_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_ab_4__13_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_5__12_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_5__12_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_5_11 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_5__11_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_4__11_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_4__12_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_5__11_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_5__11_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_5_10 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_5__10_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_4__10_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_4__11_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_5__10_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_5__10_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_5_9 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_5__9_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_4__9_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_4__10_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_5__9_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_5__9_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_5_8 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_5__8_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_4__8_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_4__9_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_5__8_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_5__8_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_5_7 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_5__7_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_4__7_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_4__8_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_5__7_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_5__7_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_5_6 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_5__6_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_4__6_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_4__7_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_5__6_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_5__6_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_5_5 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_5__5_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_4__5_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_4__6_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_5__5_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_5__5_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_5_4 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_5__4_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_4__4_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_4__5_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_5__4_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_5__4_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_5_3 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_5__3_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_4__3_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_4__4_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_5__3_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_5__3_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_5_2 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_5__2_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_4__2_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_4__3_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_5__2_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_5__2_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_5_1 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_5__1_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_4__1_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_4__2_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_5__1_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_5__1_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S1_5_0 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_5__0_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_4__0_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_4__1_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_5__0_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_A1_3_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S3_6_12 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_6__12_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_5__12_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_ab_5__13_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_6__12_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_6__12_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_6_11 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_6__11_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_5__11_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_5__12_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_6__11_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_6__11_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_6_10 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_6__10_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_5__10_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_5__11_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_6__10_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_6__10_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_6_9 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_6__9_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_5__9_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_5__10_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_6__9_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_6__9_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_6_8 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_6__8_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_5__8_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_5__9_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_6__8_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_6__8_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_6_7 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_6__7_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_5__7_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_5__8_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_6__7_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_6__7_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_6_6 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_6__6_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_5__6_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_5__7_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_6__6_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_6__6_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_6_5 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_6__5_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_5__5_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_5__6_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_6__5_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_6__5_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_6_4 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_6__4_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_5__4_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_5__5_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_6__4_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_6__4_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_6_3 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_6__3_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_5__3_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_5__4_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_6__3_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_6__3_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_6_2 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_6__2_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_5__2_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_5__3_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_6__2_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_6__2_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_6_1 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_6__1_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_5__1_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_5__2_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_6__1_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_6__1_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S1_6_0 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_6__0_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_5__0_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_5__1_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_6__0_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_A1_4_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S3_7_12 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_7__12_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_6__12_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_ab_6__13_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_7__12_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_7__12_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_7_11 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_7__11_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_6__11_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_6__12_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_7__11_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_7__11_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_7_10 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_7__10_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_6__10_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_6__11_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_7__10_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_7__10_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_7_9 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_7__9_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_6__9_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_6__10_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_7__9_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_7__9_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_7_8 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_7__8_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_6__8_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_6__9_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_7__8_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_7__8_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_7_7 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_7__7_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_6__7_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_6__8_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_7__7_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_7__7_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_7_6 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_7__6_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_6__6_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_6__7_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_7__6_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_7__6_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_7_5 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_7__5_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_6__5_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_6__6_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_7__5_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_7__5_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_7_4 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_7__4_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_6__4_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_6__5_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_7__4_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_7__4_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_7_3 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_7__3_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_6__3_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_6__4_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_7__3_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_7__3_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_7_2 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_7__2_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_6__2_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_6__3_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_7__2_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_7__2_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_7_1 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_7__1_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_6__1_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_6__2_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_7__1_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_7__1_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S1_7_0 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_7__0_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_6__0_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_6__1_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_7__0_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_A1_5_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S3_8_12 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_8__12_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_7__12_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_ab_7__13_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_8__12_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_8__12_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_8_11 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_8__11_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_7__11_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_7__12_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_8__11_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_8__11_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_8_10 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_8__10_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_7__10_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_7__11_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_8__10_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_8__10_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_8_9 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_8__9_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_7__9_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_7__10_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_8__9_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_8__9_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_8_8 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_8__8_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_7__8_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_7__9_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_8__8_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_8__8_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_8_7 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_8__7_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_7__7_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_7__8_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_8__7_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_8__7_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_8_6 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_8__6_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_7__6_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_7__7_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_8__6_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_8__6_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_8_5 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_8__5_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_7__5_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_7__6_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_8__5_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_8__5_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_8_4 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_8__4_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_7__4_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_7__5_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_8__4_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_8__4_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_8_3 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_8__3_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_7__3_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_7__4_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_8__3_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_8__3_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_8_2 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_8__2_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_7__2_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_7__3_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_8__2_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_8__2_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_8_1 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_8__1_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_7__1_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_7__2_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_8__1_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_8__1_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S1_8_0 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_8__0_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_7__0_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_7__1_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_8__0_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_A1_6_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S3_9_12 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_9__12_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_8__12_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_ab_8__13_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_9__12_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_9__12_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_9_11 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_9__11_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_8__11_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_8__12_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_9__11_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_9__11_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_9_10 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_9__10_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_8__10_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_8__11_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_9__10_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_9__10_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_9_9 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_9__9_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_8__9_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_8__10_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_9__9_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_9__9_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_9_8 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_9__8_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_8__8_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_8__9_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_9__8_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_9__8_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_9_7 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_9__7_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_8__7_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_8__8_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_9__7_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_9__7_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_9_6 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_9__6_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_8__6_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_8__7_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_9__6_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_9__6_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_9_5 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_9__5_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_8__5_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_8__6_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_9__5_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_9__5_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_9_4 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_9__4_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_8__4_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_8__5_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_9__4_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_9__4_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_9_3 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_9__3_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_8__3_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_8__4_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_9__3_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_9__3_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_9_2 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_9__2_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_8__2_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_8__3_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_9__2_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_9__2_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_9_1 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_9__1_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_8__1_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_8__2_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_9__1_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_9__1_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S1_9_0 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_9__0_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_8__0_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_8__1_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_9__0_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_A1_7_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S3_10_12 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_10__12_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_9__12_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_ab_9__13_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_10__12_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_10__12_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_10_11 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_10__11_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_9__11_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_9__12_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_10__11_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_10__11_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_10_10 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_10__10_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_9__10_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_9__11_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_10__10_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_10__10_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_10_9 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_10__9_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_9__9_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_9__10_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_10__9_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_10__9_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_10_8 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_10__8_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_9__8_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_9__9_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_10__8_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_10__8_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_10_7 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_10__7_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_9__7_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_9__8_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_10__7_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_10__7_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_10_6 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_10__6_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_9__6_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_9__7_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_10__6_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_10__6_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_10_5 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_10__5_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_9__5_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_9__6_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_10__5_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_10__5_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_10_4 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_10__4_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_9__4_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_9__5_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_10__4_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_10__4_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_10_3 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_10__3_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_9__3_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_9__4_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_10__3_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_10__3_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_10_2 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_10__2_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_9__2_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_9__3_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_10__2_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_10__2_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_10_1 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_10__1_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_9__1_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_9__2_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_10__1_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_10__1_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S1_10_0 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_10__0_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_9__0_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_9__1_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_10__0_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_A1_8_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S3_11_12 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_11__12_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_10__12_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_ab_10__13_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_11__12_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_11__12_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_11_11 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_11__11_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_10__11_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_10__12_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_11__11_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_11__11_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_11_10 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_11__10_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_10__10_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_10__11_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_11__10_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_11__10_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_11_9 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_11__9_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_10__9_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_10__10_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_11__9_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_11__9_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_11_8 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_11__8_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_10__8_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_10__9_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_11__8_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_11__8_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_11_7 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_11__7_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_10__7_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_10__8_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_11__7_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_11__7_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_11_6 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_11__6_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_10__6_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_10__7_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_11__6_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_11__6_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_11_5 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_11__5_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_10__5_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_10__6_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_11__5_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_11__5_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_11_4 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_11__4_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_10__4_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_10__5_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_11__4_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_11__4_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_11_3 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_11__3_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_10__3_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_10__4_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_11__3_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_11__3_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_11_2 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_11__2_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_10__2_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_10__3_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_11__2_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_11__2_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_11_1 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_11__1_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_10__1_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_10__2_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_11__1_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_11__1_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S1_11_0 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_11__0_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_10__0_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_10__1_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_11__0_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_A1_9_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S3_12_12 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_12__12_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_11__12_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_ab_11__13_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_12__12_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_12__12_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_12_11 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_12__11_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_11__11_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_11__12_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_12__11_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_12__11_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_12_10 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_12__10_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_11__10_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_11__11_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_12__10_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_12__10_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_12_9 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_12__9_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_11__9_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_11__10_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_12__9_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_12__9_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_12_8 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_12__8_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_11__8_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_11__9_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_12__8_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_12__8_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_12_7 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_12__7_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_11__7_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_11__8_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_12__7_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_12__7_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_12_6 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_12__6_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_11__6_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_11__7_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_12__6_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_12__6_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_12_5 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_12__5_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_11__5_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_11__6_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_12__5_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_12__5_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_12_4 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_12__4_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_11__4_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_11__5_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_12__4_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_12__4_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_12_3 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_12__3_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_11__3_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_11__4_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_12__3_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_12__3_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_12_2 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_12__2_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_11__2_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_11__3_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_12__2_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_12__2_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S2_12_1 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_12__1_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_11__1_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_11__2_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_12__1_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_12__1_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S1_12_0 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_12__0_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_11__0_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_11__1_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_12__0_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_A1_10_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S14_13 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_n86), .B(
        my_filter_adder_mult_2_multiplication_mult_21_n100), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_ab_13__13_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_13__13_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_13__13_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S5_12 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_13__12_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_12__12_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_ab_12__13_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_13__12_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_13__12_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S4_11 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_13__11_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_12__11_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_12__12_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_13__11_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_13__11_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S4_10 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_13__10_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_12__10_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_12__11_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_13__10_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_13__10_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S4_9 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_13__9_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_12__9_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_12__10_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_13__9_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_13__9_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S4_8 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_13__8_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_12__8_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_12__9_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_13__8_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_13__8_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S4_7 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_13__7_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_12__7_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_12__8_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_13__7_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_13__7_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S4_6 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_13__6_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_12__6_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_12__7_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_13__6_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_13__6_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S4_5 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_13__5_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_12__5_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_12__6_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_13__5_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_13__5_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S4_4 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_13__4_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_12__4_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_12__5_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_13__4_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_13__4_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S4_3 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_13__3_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_12__3_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_12__4_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_13__3_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_13__3_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S4_2 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_13__2_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_12__2_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_12__3_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_13__2_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_13__2_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S4_1 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_13__1_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_12__1_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_12__2_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_13__1_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_13__1_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S4_0 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_ab_13__0_), .B(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_12__0_), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_12__1_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_CARRYB_13__0_), .S(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_13__0_) );
  FA_X1 my_filter_adder_mult_2_multiplication_mult_21_S14_13_0 ( .A(
        my_filter_q_reg_chain_3__13_), .B(my_filter_q_reg_coeff[111]), .CI(
        my_filter_adder_mult_2_multiplication_mult_21_SUMB_13__0_), .CO(
        my_filter_adder_mult_2_multiplication_mult_21_A2_12_), .S(
        my_filter_adder_mult_2_res_mult[0]) );
  NAND2_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U72 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_A2_12_), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n28), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n56) );
  OAI21_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U71 ( .B1(
        my_filter_adder_mult_2_multiplication_mult_21_A2_12_), .B2(
        my_filter_adder_mult_2_multiplication_mult_21_n28), .A(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n56), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n59) );
  INV_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U70 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n59), .ZN(
        my_filter_adder_mult_2_res_mult[1]) );
  AND2_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U69 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n50), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n47), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n20) );
  AND2_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U68 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n49), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n41), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n28) );
  AND2_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U66 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n48), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n39), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n36) );
  NAND2_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U65 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n45), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n42), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n17) );
  NAND2_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U64 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n44), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n40), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n25) );
  NAND2_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U63 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n43), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n38), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n33) );
  NAND2_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U61 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n46), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n34), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n41) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U60 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n45), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n42), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n15) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U59 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n44), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n40), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n23) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U58 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n43), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n38), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n31) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U56 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n46), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n34), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n39) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U55 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n50), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n47), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n21) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U54 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n49), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n41), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n29) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U53 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n48), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n39), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n37) );
  AND2_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U51 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n31), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n30), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n44) );
  AND2_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U50 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n37), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n29), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n52) );
  NAND2_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U49 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n36), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n33), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n49) );
  NAND2_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U48 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n35), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n32), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n57) );
  INV_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U46 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n55), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n60) );
  NAND2_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U45 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n60), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n57), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n58) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U44 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n36), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n33), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n47) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U43 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n35), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n32), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n55) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U41 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n31), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n30), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n45) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U40 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_n37), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_n29), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n53) );
  OAI21_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U39 ( .B1(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n55), .B2(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n56), .A(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n57), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n51) );
  OAI21_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U38 ( .B1(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n15), .B2(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n16), .A(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n17), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n13) );
  INV_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U36 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n15), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n62) );
  NAND2_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U35 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n62), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n17), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n18) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U34 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n20), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n21), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n22) );
  INV_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U33 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n23), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n64) );
  NAND2_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U31 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n64), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n25), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n26) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U30 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n28), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n29), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n30) );
  INV_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U29 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n31), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n70) );
  NAND2_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U28 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n70), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n33), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n34) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U26 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n36), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n37), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n38) );
  INV_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U25 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n39), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n68) );
  NAND2_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U24 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n68), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n41), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n42) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U23 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n44), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n45), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n46) );
  INV_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U21 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n47), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n66) );
  NAND2_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U20 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n66), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n49), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n50) );
  NOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U19 ( .A1(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n52), .A2(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n53), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n54) );
  OAI21_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U18 ( .B1(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n23), .B2(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n24), .A(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n25), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n19) );
  OAI21_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U16 ( .B1(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n31), .B2(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n32), .A(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n33), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n27) );
  OAI21_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U13 ( .B1(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n39), .B2(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n40), .A(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n41), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n35) );
  OAI21_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U12 ( .B1(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n47), .B2(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n48), .A(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n49), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n43) );
  INV_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U11 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n21), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n63) );
  AOI21_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U10 ( .B1(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n63), .B2(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n19), .A(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n20), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n16) );
  INV_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U9 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n29), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n71) );
  AOI21_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U8 ( .B1(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n71), .B2(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n27), .A(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n28), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n24) );
  INV_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U7 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n37), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n69) );
  AOI21_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U6 ( .B1(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n69), .B2(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n35), .A(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n36), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n32) );
  INV_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U5 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n45), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n67) );
  AOI21_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U4 ( .B1(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n67), .B2(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n43), .A(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n44), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n40) );
  INV_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U3 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n53), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n65) );
  AOI21_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U2 ( .B1(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n65), .B2(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n51), .A(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n52), .ZN(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n48) );
  XOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U67 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n56), .B(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n58), .Z(
        my_filter_adder_mult_2_res_mult[2]) );
  XOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U62 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n51), .B(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n54), .Z(
        my_filter_adder_mult_2_res_mult[3]) );
  XOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U57 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n50), .B(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n48), .Z(
        my_filter_adder_mult_2_res_mult[4]) );
  XOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U52 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n43), .B(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n46), .Z(
        my_filter_adder_mult_2_res_mult[5]) );
  XOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U47 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n42), .B(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n40), .Z(
        my_filter_adder_mult_2_res_mult[6]) );
  XOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U42 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n35), .B(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n38), .Z(
        my_filter_adder_mult_2_res_mult[7]) );
  XOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U37 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n34), .B(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n32), .Z(
        my_filter_adder_mult_2_res_mult[8]) );
  XOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U32 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n27), .B(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n30), .Z(
        my_filter_adder_mult_2_res_mult[9]) );
  XOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U27 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n26), .B(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n24), .Z(
        my_filter_adder_mult_2_res_mult[10]) );
  XOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U22 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n19), .B(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n22), .Z(
        my_filter_adder_mult_2_res_mult[11]) );
  XOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U17 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n18), .B(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n16), .Z(
        my_filter_adder_mult_2_res_mult[12]) );
  XOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U15 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_n52), .B(
        my_filter_adder_mult_2_multiplication_mult_21_n51), .Z(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n14) );
  XOR2_X1 my_filter_adder_mult_2_multiplication_mult_21_FS_1_U14 ( .A(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n13), .B(
        my_filter_adder_mult_2_multiplication_mult_21_FS_1_n14), .Z(
        my_filter_adder_mult_2_res_mult[13]) );
  AND2_X1 my_filter_adder_mult_2_addition_add_19_U1 ( .A1(
        my_filter_data_sum[112]), .A2(my_filter_adder_mult_2_res_mult[0]), 
        .ZN(my_filter_adder_mult_2_addition_add_19_n1) );
  XOR2_X1 my_filter_adder_mult_2_addition_add_19_U2 ( .A(
        my_filter_data_sum[112]), .B(my_filter_adder_mult_2_res_mult[0]), .Z(
        my_filter_data_sum[98]) );
  FA_X1 my_filter_adder_mult_2_addition_add_19_U1_1 ( .A(
        my_filter_adder_mult_2_res_mult[1]), .B(my_filter_data_sum[113]), .CI(
        my_filter_adder_mult_2_addition_add_19_n1), .CO(
        my_filter_adder_mult_2_addition_add_19_carry[2]), .S(
        my_filter_data_sum[99]) );
  FA_X1 my_filter_adder_mult_2_addition_add_19_U1_2 ( .A(
        my_filter_adder_mult_2_res_mult[2]), .B(my_filter_data_sum[114]), .CI(
        my_filter_adder_mult_2_addition_add_19_carry[2]), .CO(
        my_filter_adder_mult_2_addition_add_19_carry[3]), .S(
        my_filter_data_sum[100]) );
  FA_X1 my_filter_adder_mult_2_addition_add_19_U1_3 ( .A(
        my_filter_adder_mult_2_res_mult[3]), .B(my_filter_data_sum[115]), .CI(
        my_filter_adder_mult_2_addition_add_19_carry[3]), .CO(
        my_filter_adder_mult_2_addition_add_19_carry[4]), .S(
        my_filter_data_sum[101]) );
  FA_X1 my_filter_adder_mult_2_addition_add_19_U1_4 ( .A(
        my_filter_adder_mult_2_res_mult[4]), .B(my_filter_data_sum[116]), .CI(
        my_filter_adder_mult_2_addition_add_19_carry[4]), .CO(
        my_filter_adder_mult_2_addition_add_19_carry[5]), .S(
        my_filter_data_sum[102]) );
  FA_X1 my_filter_adder_mult_2_addition_add_19_U1_5 ( .A(
        my_filter_adder_mult_2_res_mult[5]), .B(my_filter_data_sum[117]), .CI(
        my_filter_adder_mult_2_addition_add_19_carry[5]), .CO(
        my_filter_adder_mult_2_addition_add_19_carry[6]), .S(
        my_filter_data_sum[103]) );
  FA_X1 my_filter_adder_mult_2_addition_add_19_U1_6 ( .A(
        my_filter_adder_mult_2_res_mult[6]), .B(my_filter_data_sum[118]), .CI(
        my_filter_adder_mult_2_addition_add_19_carry[6]), .CO(
        my_filter_adder_mult_2_addition_add_19_carry[7]), .S(
        my_filter_data_sum[104]) );
  FA_X1 my_filter_adder_mult_2_addition_add_19_U1_7 ( .A(
        my_filter_adder_mult_2_res_mult[7]), .B(my_filter_data_sum[119]), .CI(
        my_filter_adder_mult_2_addition_add_19_carry[7]), .CO(
        my_filter_adder_mult_2_addition_add_19_carry[8]), .S(
        my_filter_data_sum[105]) );
  FA_X1 my_filter_adder_mult_2_addition_add_19_U1_8 ( .A(
        my_filter_adder_mult_2_res_mult[8]), .B(my_filter_data_sum[120]), .CI(
        my_filter_adder_mult_2_addition_add_19_carry[8]), .CO(
        my_filter_adder_mult_2_addition_add_19_carry[9]), .S(
        my_filter_data_sum[106]) );
  FA_X1 my_filter_adder_mult_2_addition_add_19_U1_9 ( .A(
        my_filter_adder_mult_2_res_mult[9]), .B(my_filter_data_sum[121]), .CI(
        my_filter_adder_mult_2_addition_add_19_carry[9]), .CO(
        my_filter_adder_mult_2_addition_add_19_carry[10]), .S(
        my_filter_data_sum[107]) );
  FA_X1 my_filter_adder_mult_2_addition_add_19_U1_10 ( .A(
        my_filter_adder_mult_2_res_mult[10]), .B(my_filter_data_sum[122]), 
        .CI(my_filter_adder_mult_2_addition_add_19_carry[10]), .CO(
        my_filter_adder_mult_2_addition_add_19_carry[11]), .S(
        my_filter_data_sum[108]) );
  FA_X1 my_filter_adder_mult_2_addition_add_19_U1_11 ( .A(
        my_filter_adder_mult_2_res_mult[11]), .B(my_filter_data_sum[123]), 
        .CI(my_filter_adder_mult_2_addition_add_19_carry[11]), .CO(
        my_filter_adder_mult_2_addition_add_19_carry[12]), .S(
        my_filter_data_sum[109]) );
  FA_X1 my_filter_adder_mult_2_addition_add_19_U1_12 ( .A(
        my_filter_adder_mult_2_res_mult[12]), .B(my_filter_data_sum[124]), 
        .CI(my_filter_adder_mult_2_addition_add_19_carry[12]), .CO(
        my_filter_adder_mult_2_addition_add_19_carry[13]), .S(
        my_filter_data_sum[110]) );
  FA_X1 my_filter_adder_mult_2_addition_add_19_U1_13 ( .A(
        my_filter_adder_mult_2_res_mult[13]), .B(my_filter_data_sum[125]), 
        .CI(my_filter_adder_mult_2_addition_add_19_carry[13]), .S(
        my_filter_data_sum[111]) );
  INV_X1 my_filter_adder_mult_3_multiplication_mult_21_U276 ( .A(
        my_filter_q_reg_chain_4__13_), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_n86) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U275 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_12__12_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U274 ( .A1(
        my_filter_q_reg_chain_4__11_), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_11__13_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U273 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_11__12_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U272 ( .A1(
        my_filter_q_reg_chain_4__10_), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_10__13_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U271 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_10__12_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U270 ( .A1(
        my_filter_q_reg_chain_4__9_), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_9__13_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U269 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n101), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_9__12_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U268 ( .A1(
        my_filter_q_reg_chain_4__8_), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_8__13_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U267 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_8__12_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U266 ( .A1(
        my_filter_q_reg_chain_4__7_), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_7__13_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U265 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_7__12_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U264 ( .A1(
        my_filter_q_reg_chain_4__6_), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_6__13_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U263 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_6__12_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U262 ( .A1(
        my_filter_q_reg_chain_4__5_), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_5__13_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U261 ( .A1(
        my_filter_q_reg_coeff[95]), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_13__11_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U260 ( .A1(
        my_filter_q_reg_coeff[94]), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_13__10_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U259 ( .A1(
        my_filter_q_reg_coeff[92]), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_13__8_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U258 ( .A1(
        my_filter_q_reg_coeff[93]), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_13__9_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U257 ( .A1(
        my_filter_q_reg_coeff[90]), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_13__6_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U256 ( .A1(
        my_filter_q_reg_coeff[91]), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_13__7_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U255 ( .A1(
        my_filter_q_reg_coeff[89]), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_13__5_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U254 ( .A1(
        my_filter_q_reg_coeff[96]), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_13__12_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U253 ( .A1(
        my_filter_q_reg_chain_4__12_), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_12__13_) );
  INV_X1 my_filter_adder_mult_3_multiplication_mult_21_U252 ( .A(
        my_filter_q_reg_chain_4__9_), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_n90) );
  INV_X1 my_filter_adder_mult_3_multiplication_mult_21_U251 ( .A(
        my_filter_q_reg_chain_4__12_), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_n87) );
  INV_X1 my_filter_adder_mult_3_multiplication_mult_21_U250 ( .A(
        my_filter_q_reg_chain_4__11_), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_n88) );
  INV_X1 my_filter_adder_mult_3_multiplication_mult_21_U249 ( .A(
        my_filter_q_reg_chain_4__10_), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_n89) );
  INV_X1 my_filter_adder_mult_3_multiplication_mult_21_U248 ( .A(
        my_filter_q_reg_chain_4__8_), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_n91) );
  INV_X1 my_filter_adder_mult_3_multiplication_mult_21_U247 ( .A(
        my_filter_q_reg_chain_4__7_), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_n92) );
  INV_X1 my_filter_adder_mult_3_multiplication_mult_21_U246 ( .A(
        my_filter_q_reg_chain_4__6_), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_n93) );
  INV_X1 my_filter_adder_mult_3_multiplication_mult_21_U245 ( .A(
        my_filter_q_reg_chain_4__5_), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_n94) );
  AND2_X1 my_filter_adder_mult_3_multiplication_mult_21_U244 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_ab_0__13_), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_ab_1__12_), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_n15) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U243 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_2__12_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U242 ( .A1(
        my_filter_q_reg_chain_4__1_), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_1__13_) );
  AND3_X1 my_filter_adder_mult_3_multiplication_mult_21_U241 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_ab_1__1_), .A2(
        my_filter_q_reg_coeff[84]), .A3(my_filter_q_reg_chain_4__0_), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_1__0_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U240 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_12__0_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U239 ( .A1(
        my_filter_q_reg_coeff[84]), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_13__0_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U238 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_5__12_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U237 ( .A1(
        my_filter_q_reg_chain_4__4_), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_4__13_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U236 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_4__12_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U235 ( .A1(
        my_filter_q_reg_chain_4__3_), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_3__13_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U234 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_3__12_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U233 ( .A1(
        my_filter_q_reg_chain_4__2_), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_2__13_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U232 ( .A1(
        my_filter_q_reg_coeff[88]), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_13__4_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U231 ( .A1(
        my_filter_q_reg_coeff[85]), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_13__1_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U230 ( .A1(
        my_filter_q_reg_coeff[86]), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_13__2_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U229 ( .A1(
        my_filter_q_reg_coeff[87]), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_13__3_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U228 ( .A1(
        my_filter_q_reg_chain_4__0_), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_0__13_) );
  INV_X1 my_filter_adder_mult_3_multiplication_mult_21_U227 ( .A(
        my_filter_q_reg_coeff[97]), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_n100) );
  INV_X1 my_filter_adder_mult_3_multiplication_mult_21_U226 ( .A(
        my_filter_q_reg_coeff[84]), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_n113) );
  INV_X1 my_filter_adder_mult_3_multiplication_mult_21_U225 ( .A(
        my_filter_q_reg_chain_4__0_), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_n99) );
  INV_X1 my_filter_adder_mult_3_multiplication_mult_21_U224 ( .A(
        my_filter_q_reg_coeff[85]), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_n112) );
  INV_X1 my_filter_adder_mult_3_multiplication_mult_21_U223 ( .A(
        my_filter_q_reg_chain_4__1_), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_n98) );
  INV_X1 my_filter_adder_mult_3_multiplication_mult_21_U222 ( .A(
        my_filter_q_reg_coeff[96]), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_n101) );
  INV_X1 my_filter_adder_mult_3_multiplication_mult_21_U221 ( .A(
        my_filter_q_reg_coeff[94]), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_n103) );
  INV_X1 my_filter_adder_mult_3_multiplication_mult_21_U220 ( .A(
        my_filter_q_reg_coeff[95]), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_n102) );
  INV_X1 my_filter_adder_mult_3_multiplication_mult_21_U219 ( .A(
        my_filter_q_reg_coeff[92]), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_n105) );
  INV_X1 my_filter_adder_mult_3_multiplication_mult_21_U218 ( .A(
        my_filter_q_reg_coeff[93]), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_n104) );
  INV_X1 my_filter_adder_mult_3_multiplication_mult_21_U217 ( .A(
        my_filter_q_reg_coeff[89]), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_n108) );
  INV_X1 my_filter_adder_mult_3_multiplication_mult_21_U216 ( .A(
        my_filter_q_reg_coeff[90]), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_n107) );
  INV_X1 my_filter_adder_mult_3_multiplication_mult_21_U215 ( .A(
        my_filter_q_reg_coeff[91]), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_n106) );
  INV_X1 my_filter_adder_mult_3_multiplication_mult_21_U214 ( .A(
        my_filter_q_reg_coeff[86]), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_n111) );
  INV_X1 my_filter_adder_mult_3_multiplication_mult_21_U213 ( .A(
        my_filter_q_reg_coeff[87]), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_n110) );
  INV_X1 my_filter_adder_mult_3_multiplication_mult_21_U212 ( .A(
        my_filter_q_reg_coeff[88]), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_n109) );
  INV_X1 my_filter_adder_mult_3_multiplication_mult_21_U211 ( .A(
        my_filter_q_reg_chain_4__4_), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_n95) );
  INV_X1 my_filter_adder_mult_3_multiplication_mult_21_U210 ( .A(
        my_filter_q_reg_chain_4__2_), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_n97) );
  INV_X1 my_filter_adder_mult_3_multiplication_mult_21_U209 ( .A(
        my_filter_q_reg_chain_4__3_), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_n96) );
  AND2_X1 my_filter_adder_mult_3_multiplication_mult_21_U208 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_13__12_), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_13__13_), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_n3) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U207 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n100), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_13__13_) );
  AND2_X1 my_filter_adder_mult_3_multiplication_mult_21_U206 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_13__9_), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_13__10_), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_n51) );
  AND2_X1 my_filter_adder_mult_3_multiplication_mult_21_U205 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_13__7_), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_13__8_), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_n50) );
  AND2_X1 my_filter_adder_mult_3_multiplication_mult_21_U204 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_13__5_), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_13__6_), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_n49) );
  AND2_X1 my_filter_adder_mult_3_multiplication_mult_21_U203 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_13__3_), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_13__4_), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_n42) );
  AND2_X1 my_filter_adder_mult_3_multiplication_mult_21_U202 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_13__10_), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_13__11_), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_n44) );
  AND2_X1 my_filter_adder_mult_3_multiplication_mult_21_U201 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_13__8_), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_13__9_), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_n43) );
  AND2_X1 my_filter_adder_mult_3_multiplication_mult_21_U200 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_13__6_), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_13__7_), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_n47) );
  AND2_X1 my_filter_adder_mult_3_multiplication_mult_21_U199 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_13__4_), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_13__5_), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_n46) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U198 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_12__11_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U197 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_12__9_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U196 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_12__10_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U195 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_11__10_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U194 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_11__11_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U193 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_12__7_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U192 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_12__8_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U191 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_10__11_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U190 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_11__8_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U189 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_11__9_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U188 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_12__6_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U187 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_10__9_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U186 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_10__10_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U185 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_11__7_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U184 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n103), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_9__10_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U183 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n102), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_9__11_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U182 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_10__8_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U181 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_8__11_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U180 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n104), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_9__9_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U179 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_8__10_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U178 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_7__11_) );
  AND2_X1 my_filter_adder_mult_3_multiplication_mult_21_U177 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_13__11_), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_13__12_), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_n52) );
  AND2_X1 my_filter_adder_mult_3_multiplication_mult_21_U176 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_13__1_), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_13__2_), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_n35) );
  AND2_X1 my_filter_adder_mult_3_multiplication_mult_21_U175 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_13__2_), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_13__3_), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_n34) );
  AND2_X1 my_filter_adder_mult_3_multiplication_mult_21_U174 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_13__0_), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_13__1_), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_n33) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U173 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_12__1_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U172 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_10__0_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U171 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_11__0_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U170 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_11__1_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U169 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_10__1_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U168 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_8__0_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U167 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n113), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_9__0_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U166 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n112), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_9__1_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U165 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n110), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_9__3_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U164 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_8__1_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U163 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_8__3_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U162 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_6__0_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U161 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_7__0_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U160 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_7__1_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U159 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_7__3_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U158 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_7__4_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U157 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_7__5_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U156 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_6__1_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U155 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_6__3_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U154 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_6__5_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U153 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_4__0_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U152 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_5__0_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U151 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_5__1_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U150 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_5__3_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U149 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_5__4_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U148 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_5__5_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U147 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_5__6_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U146 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_4__1_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U145 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_4__3_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U144 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_4__5_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U143 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_2__0_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U142 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_3__0_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U141 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_3__1_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U140 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_3__3_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U139 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_3__4_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U138 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_3__5_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U137 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_3__6_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U136 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_3__7_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U135 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_12__5_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U134 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_11__6_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U133 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_12__2_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U132 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_12__3_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U131 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_12__4_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U130 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_10__7_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U129 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_11__3_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U128 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_11__4_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U127 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_11__5_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U126 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n105), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_9__8_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U125 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_10__4_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U124 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_10__5_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U123 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_10__6_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U122 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_8__9_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U121 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_11__2_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U120 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n108), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_9__5_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U119 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n107), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_9__6_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U118 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n106), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_9__7_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U117 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_7__10_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U116 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_10__2_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U115 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_10__3_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U114 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_8__6_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U113 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_8__7_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U112 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_8__8_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U111 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_6__11_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U110 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n111), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_9__2_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U109 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n109), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_9__4_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U108 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_7__7_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U107 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_7__8_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U106 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_7__9_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U105 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_8__2_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U104 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_8__4_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U103 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_8__5_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U102 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_6__8_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U101 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_6__9_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U100 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_6__10_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U99 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_7__2_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U98 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_7__6_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U97 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_5__9_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U96 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_5__10_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U95 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_5__11_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U94 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_6__2_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U93 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_6__4_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U92 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_6__6_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U91 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_6__7_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U90 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_4__10_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U89 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_4__11_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U88 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_5__2_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U87 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_5__7_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U86 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_5__8_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U85 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_3__11_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U84 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_4__2_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U83 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_4__4_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U82 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_4__6_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U81 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_4__7_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U80 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_4__8_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U79 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_4__9_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U78 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_3__2_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U77 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_3__8_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U76 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_3__9_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U75 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_3__10_) );
  AND2_X1 my_filter_adder_mult_3_multiplication_mult_21_U74 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_ab_0__2_), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_ab_1__1_), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_n14) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U73 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_2__1_) );
  AND2_X1 my_filter_adder_mult_3_multiplication_mult_21_U72 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_ab_0__3_), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_ab_1__2_), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_n13) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U71 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_2__2_) );
  AND2_X1 my_filter_adder_mult_3_multiplication_mult_21_U70 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_ab_0__4_), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_ab_1__3_), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_n12) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U69 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_2__3_) );
  AND2_X1 my_filter_adder_mult_3_multiplication_mult_21_U68 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_ab_0__5_), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_ab_1__4_), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_n11) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U67 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_2__4_) );
  AND2_X1 my_filter_adder_mult_3_multiplication_mult_21_U66 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_ab_0__6_), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_ab_1__5_), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_n10) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U65 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_2__5_) );
  AND2_X1 my_filter_adder_mult_3_multiplication_mult_21_U64 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_ab_0__7_), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_ab_1__6_), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_n9) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U63 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_2__6_) );
  AND2_X1 my_filter_adder_mult_3_multiplication_mult_21_U62 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_ab_0__8_), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_ab_1__7_), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_n8) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U61 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_2__7_) );
  AND2_X1 my_filter_adder_mult_3_multiplication_mult_21_U60 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_ab_0__9_), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_ab_1__8_), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_n7) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U59 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_2__8_) );
  AND2_X1 my_filter_adder_mult_3_multiplication_mult_21_U58 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_ab_0__10_), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_ab_1__9_), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_n6) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U57 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_2__9_) );
  AND2_X1 my_filter_adder_mult_3_multiplication_mult_21_U56 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_ab_0__11_), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_ab_1__10_), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_n5) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U55 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_2__10_) );
  AND2_X1 my_filter_adder_mult_3_multiplication_mult_21_U54 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_ab_0__12_), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_ab_1__11_), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_n4) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U52 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_2__11_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U51 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_1__12_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U50 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_1__2_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U49 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_1__3_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U47 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_1__4_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U46 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_1__5_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U44 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_1__6_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U43 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_1__7_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U42 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_1__8_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U35 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_1__9_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U34 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_1__10_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U33 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_1__11_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U14 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_0__2_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U13 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_0__3_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U12 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_0__4_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U11 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_0__5_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U10 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_0__6_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U9 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_0__7_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U8 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_0__8_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U7 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_0__9_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U6 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_0__10_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U5 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_0__11_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U4 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_0__12_) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U3 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n98), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n112), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_ab_1__1_) );
  INV_X1 my_filter_adder_mult_3_multiplication_mult_21_U2 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_13__13_), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_n85) );
  XOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U48 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_13__10_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_13__11_), .Z(
        my_filter_adder_mult_3_multiplication_mult_21_n48) );
  XOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U45 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_13__5_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_13__6_), .Z(
        my_filter_adder_mult_3_multiplication_mult_21_n45) );
  XOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U41 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_13__11_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_13__12_), .Z(
        my_filter_adder_mult_3_multiplication_mult_21_n41) );
  XOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U40 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_13__8_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_13__9_), .Z(
        my_filter_adder_mult_3_multiplication_mult_21_n40) );
  XOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U39 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_13__9_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_13__10_), .Z(
        my_filter_adder_mult_3_multiplication_mult_21_n39) );
  XOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U38 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_13__6_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_13__7_), .Z(
        my_filter_adder_mult_3_multiplication_mult_21_n38) );
  XOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U37 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_13__7_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_13__8_), .Z(
        my_filter_adder_mult_3_multiplication_mult_21_n37) );
  XOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U36 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_13__4_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_13__5_), .Z(
        my_filter_adder_mult_3_multiplication_mult_21_n36) );
  XOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U32 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_13__3_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_13__4_), .Z(
        my_filter_adder_mult_3_multiplication_mult_21_n32) );
  XOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U31 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_13__1_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_13__2_), .Z(
        my_filter_adder_mult_3_multiplication_mult_21_n31) );
  XOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U30 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_13__2_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_13__3_), .Z(
        my_filter_adder_mult_3_multiplication_mult_21_n30) );
  XOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U29 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_13__0_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_13__1_), .Z(
        my_filter_adder_mult_3_multiplication_mult_21_n29) );
  XOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U27 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_1__1_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_ab_0__2_), .Z(
        my_filter_adder_mult_3_multiplication_mult_21_n28) );
  XOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U26 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_13__12_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_13__13_), .Z(
        my_filter_adder_mult_3_multiplication_mult_21_n27) );
  XOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U25 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_1__12_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_ab_0__13_), .Z(
        my_filter_adder_mult_3_multiplication_mult_21_n26) );
  XOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U24 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_1__2_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_ab_0__3_), .Z(
        my_filter_adder_mult_3_multiplication_mult_21_n25) );
  XOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U23 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_1__3_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_ab_0__4_), .Z(
        my_filter_adder_mult_3_multiplication_mult_21_n24) );
  XOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U22 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_1__4_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_ab_0__5_), .Z(
        my_filter_adder_mult_3_multiplication_mult_21_n23) );
  XOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U21 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_1__5_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_ab_0__6_), .Z(
        my_filter_adder_mult_3_multiplication_mult_21_n22) );
  XOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U20 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_1__6_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_ab_0__7_), .Z(
        my_filter_adder_mult_3_multiplication_mult_21_n21) );
  XOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U19 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_1__7_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_ab_0__8_), .Z(
        my_filter_adder_mult_3_multiplication_mult_21_n20) );
  XOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U18 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_1__8_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_ab_0__9_), .Z(
        my_filter_adder_mult_3_multiplication_mult_21_n19) );
  XOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U17 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_1__9_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_ab_0__10_), .Z(
        my_filter_adder_mult_3_multiplication_mult_21_n18) );
  XOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U16 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_1__10_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_ab_0__11_), .Z(
        my_filter_adder_mult_3_multiplication_mult_21_n17) );
  XOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_U15 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_1__11_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_ab_0__12_), .Z(
        my_filter_adder_mult_3_multiplication_mult_21_n16) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S3_2_12 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_2__12_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_n15), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_ab_1__13_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_2__12_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_2__12_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_2_11 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_2__11_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_n4), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_n26), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_2__11_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_2__11_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_2_10 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_2__10_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_n5), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_n16), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_2__10_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_2__10_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_2_9 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_2__9_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_n6), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_n17), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_2__9_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_2__9_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_2_8 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_2__8_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_n7), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_n18), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_2__8_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_2__8_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_2_7 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_2__7_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_n8), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_n19), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_2__7_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_2__7_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_2_6 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_2__6_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_n9), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_n20), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_2__6_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_2__6_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_2_5 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_2__5_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_n10), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_n21), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_2__5_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_2__5_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_2_4 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_2__4_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_n11), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_n22), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_2__4_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_2__4_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_2_3 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_2__3_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_n12), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_n23), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_2__3_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_2__3_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_2_2 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_2__2_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_n13), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_n24), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_2__2_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_2__2_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_2_1 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_2__1_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_n14), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_n25), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_2__1_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_2__1_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S1_2_0 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_2__0_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_1__0_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_n28), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_2__0_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_A1_0_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S3_3_12 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_3__12_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_2__12_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_ab_2__13_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_3__12_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_3__12_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_3_11 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_3__11_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_2__11_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_2__12_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_3__11_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_3__11_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_3_10 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_3__10_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_2__10_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_2__11_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_3__10_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_3__10_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_3_9 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_3__9_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_2__9_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_2__10_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_3__9_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_3__9_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_3_8 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_3__8_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_2__8_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_2__9_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_3__8_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_3__8_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_3_7 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_3__7_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_2__7_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_2__8_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_3__7_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_3__7_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_3_6 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_3__6_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_2__6_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_2__7_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_3__6_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_3__6_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_3_5 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_3__5_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_2__5_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_2__6_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_3__5_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_3__5_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_3_4 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_3__4_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_2__4_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_2__5_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_3__4_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_3__4_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_3_3 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_3__3_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_2__3_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_2__4_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_3__3_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_3__3_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_3_2 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_3__2_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_2__2_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_2__3_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_3__2_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_3__2_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_3_1 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_3__1_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_2__1_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_2__2_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_3__1_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_3__1_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S1_3_0 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_3__0_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_2__0_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_2__1_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_3__0_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_A1_1_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S3_4_12 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_4__12_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_3__12_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_ab_3__13_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_4__12_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_4__12_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_4_11 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_4__11_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_3__11_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_3__12_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_4__11_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_4__11_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_4_10 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_4__10_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_3__10_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_3__11_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_4__10_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_4__10_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_4_9 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_4__9_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_3__9_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_3__10_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_4__9_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_4__9_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_4_8 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_4__8_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_3__8_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_3__9_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_4__8_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_4__8_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_4_7 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_4__7_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_3__7_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_3__8_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_4__7_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_4__7_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_4_6 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_4__6_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_3__6_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_3__7_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_4__6_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_4__6_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_4_5 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_4__5_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_3__5_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_3__6_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_4__5_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_4__5_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_4_4 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_4__4_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_3__4_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_3__5_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_4__4_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_4__4_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_4_3 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_4__3_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_3__3_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_3__4_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_4__3_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_4__3_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_4_2 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_4__2_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_3__2_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_3__3_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_4__2_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_4__2_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_4_1 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_4__1_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_3__1_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_3__2_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_4__1_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_4__1_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S1_4_0 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_4__0_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_3__0_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_3__1_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_4__0_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_A1_2_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S3_5_12 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_5__12_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_4__12_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_ab_4__13_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_5__12_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_5__12_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_5_11 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_5__11_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_4__11_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_4__12_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_5__11_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_5__11_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_5_10 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_5__10_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_4__10_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_4__11_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_5__10_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_5__10_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_5_9 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_5__9_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_4__9_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_4__10_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_5__9_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_5__9_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_5_8 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_5__8_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_4__8_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_4__9_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_5__8_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_5__8_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_5_7 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_5__7_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_4__7_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_4__8_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_5__7_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_5__7_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_5_6 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_5__6_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_4__6_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_4__7_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_5__6_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_5__6_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_5_5 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_5__5_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_4__5_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_4__6_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_5__5_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_5__5_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_5_4 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_5__4_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_4__4_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_4__5_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_5__4_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_5__4_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_5_3 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_5__3_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_4__3_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_4__4_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_5__3_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_5__3_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_5_2 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_5__2_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_4__2_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_4__3_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_5__2_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_5__2_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_5_1 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_5__1_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_4__1_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_4__2_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_5__1_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_5__1_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S1_5_0 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_5__0_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_4__0_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_4__1_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_5__0_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_A1_3_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S3_6_12 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_6__12_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_5__12_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_ab_5__13_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_6__12_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_6__12_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_6_11 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_6__11_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_5__11_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_5__12_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_6__11_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_6__11_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_6_10 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_6__10_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_5__10_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_5__11_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_6__10_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_6__10_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_6_9 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_6__9_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_5__9_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_5__10_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_6__9_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_6__9_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_6_8 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_6__8_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_5__8_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_5__9_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_6__8_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_6__8_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_6_7 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_6__7_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_5__7_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_5__8_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_6__7_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_6__7_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_6_6 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_6__6_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_5__6_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_5__7_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_6__6_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_6__6_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_6_5 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_6__5_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_5__5_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_5__6_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_6__5_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_6__5_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_6_4 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_6__4_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_5__4_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_5__5_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_6__4_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_6__4_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_6_3 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_6__3_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_5__3_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_5__4_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_6__3_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_6__3_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_6_2 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_6__2_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_5__2_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_5__3_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_6__2_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_6__2_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_6_1 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_6__1_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_5__1_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_5__2_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_6__1_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_6__1_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S1_6_0 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_6__0_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_5__0_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_5__1_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_6__0_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_A1_4_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S3_7_12 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_7__12_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_6__12_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_ab_6__13_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_7__12_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_7__12_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_7_11 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_7__11_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_6__11_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_6__12_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_7__11_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_7__11_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_7_10 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_7__10_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_6__10_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_6__11_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_7__10_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_7__10_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_7_9 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_7__9_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_6__9_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_6__10_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_7__9_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_7__9_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_7_8 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_7__8_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_6__8_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_6__9_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_7__8_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_7__8_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_7_7 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_7__7_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_6__7_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_6__8_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_7__7_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_7__7_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_7_6 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_7__6_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_6__6_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_6__7_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_7__6_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_7__6_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_7_5 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_7__5_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_6__5_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_6__6_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_7__5_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_7__5_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_7_4 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_7__4_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_6__4_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_6__5_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_7__4_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_7__4_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_7_3 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_7__3_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_6__3_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_6__4_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_7__3_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_7__3_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_7_2 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_7__2_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_6__2_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_6__3_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_7__2_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_7__2_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_7_1 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_7__1_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_6__1_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_6__2_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_7__1_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_7__1_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S1_7_0 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_7__0_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_6__0_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_6__1_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_7__0_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_A1_5_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S3_8_12 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_8__12_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_7__12_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_ab_7__13_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_8__12_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_8__12_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_8_11 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_8__11_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_7__11_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_7__12_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_8__11_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_8__11_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_8_10 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_8__10_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_7__10_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_7__11_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_8__10_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_8__10_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_8_9 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_8__9_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_7__9_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_7__10_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_8__9_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_8__9_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_8_8 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_8__8_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_7__8_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_7__9_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_8__8_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_8__8_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_8_7 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_8__7_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_7__7_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_7__8_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_8__7_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_8__7_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_8_6 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_8__6_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_7__6_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_7__7_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_8__6_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_8__6_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_8_5 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_8__5_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_7__5_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_7__6_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_8__5_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_8__5_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_8_4 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_8__4_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_7__4_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_7__5_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_8__4_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_8__4_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_8_3 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_8__3_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_7__3_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_7__4_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_8__3_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_8__3_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_8_2 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_8__2_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_7__2_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_7__3_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_8__2_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_8__2_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_8_1 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_8__1_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_7__1_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_7__2_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_8__1_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_8__1_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S1_8_0 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_8__0_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_7__0_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_7__1_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_8__0_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_A1_6_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S3_9_12 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_9__12_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_8__12_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_ab_8__13_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_9__12_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_9__12_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_9_11 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_9__11_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_8__11_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_8__12_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_9__11_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_9__11_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_9_10 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_9__10_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_8__10_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_8__11_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_9__10_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_9__10_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_9_9 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_9__9_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_8__9_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_8__10_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_9__9_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_9__9_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_9_8 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_9__8_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_8__8_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_8__9_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_9__8_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_9__8_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_9_7 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_9__7_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_8__7_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_8__8_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_9__7_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_9__7_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_9_6 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_9__6_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_8__6_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_8__7_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_9__6_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_9__6_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_9_5 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_9__5_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_8__5_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_8__6_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_9__5_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_9__5_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_9_4 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_9__4_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_8__4_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_8__5_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_9__4_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_9__4_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_9_3 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_9__3_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_8__3_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_8__4_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_9__3_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_9__3_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_9_2 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_9__2_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_8__2_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_8__3_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_9__2_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_9__2_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_9_1 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_9__1_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_8__1_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_8__2_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_9__1_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_9__1_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S1_9_0 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_9__0_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_8__0_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_8__1_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_9__0_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_A1_7_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S3_10_12 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_10__12_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_9__12_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_ab_9__13_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_10__12_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_10__12_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_10_11 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_10__11_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_9__11_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_9__12_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_10__11_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_10__11_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_10_10 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_10__10_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_9__10_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_9__11_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_10__10_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_10__10_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_10_9 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_10__9_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_9__9_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_9__10_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_10__9_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_10__9_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_10_8 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_10__8_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_9__8_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_9__9_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_10__8_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_10__8_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_10_7 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_10__7_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_9__7_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_9__8_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_10__7_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_10__7_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_10_6 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_10__6_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_9__6_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_9__7_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_10__6_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_10__6_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_10_5 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_10__5_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_9__5_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_9__6_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_10__5_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_10__5_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_10_4 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_10__4_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_9__4_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_9__5_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_10__4_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_10__4_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_10_3 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_10__3_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_9__3_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_9__4_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_10__3_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_10__3_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_10_2 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_10__2_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_9__2_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_9__3_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_10__2_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_10__2_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_10_1 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_10__1_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_9__1_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_9__2_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_10__1_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_10__1_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S1_10_0 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_10__0_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_9__0_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_9__1_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_10__0_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_A1_8_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S3_11_12 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_11__12_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_10__12_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_ab_10__13_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_11__12_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_11__12_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_11_11 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_11__11_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_10__11_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_10__12_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_11__11_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_11__11_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_11_10 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_11__10_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_10__10_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_10__11_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_11__10_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_11__10_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_11_9 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_11__9_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_10__9_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_10__10_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_11__9_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_11__9_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_11_8 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_11__8_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_10__8_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_10__9_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_11__8_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_11__8_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_11_7 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_11__7_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_10__7_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_10__8_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_11__7_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_11__7_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_11_6 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_11__6_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_10__6_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_10__7_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_11__6_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_11__6_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_11_5 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_11__5_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_10__5_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_10__6_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_11__5_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_11__5_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_11_4 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_11__4_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_10__4_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_10__5_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_11__4_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_11__4_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_11_3 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_11__3_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_10__3_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_10__4_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_11__3_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_11__3_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_11_2 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_11__2_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_10__2_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_10__3_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_11__2_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_11__2_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_11_1 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_11__1_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_10__1_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_10__2_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_11__1_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_11__1_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S1_11_0 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_11__0_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_10__0_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_10__1_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_11__0_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_A1_9_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S3_12_12 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_12__12_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_11__12_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_ab_11__13_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_12__12_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_12__12_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_12_11 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_12__11_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_11__11_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_11__12_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_12__11_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_12__11_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_12_10 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_12__10_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_11__10_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_11__11_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_12__10_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_12__10_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_12_9 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_12__9_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_11__9_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_11__10_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_12__9_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_12__9_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_12_8 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_12__8_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_11__8_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_11__9_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_12__8_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_12__8_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_12_7 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_12__7_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_11__7_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_11__8_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_12__7_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_12__7_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_12_6 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_12__6_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_11__6_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_11__7_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_12__6_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_12__6_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_12_5 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_12__5_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_11__5_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_11__6_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_12__5_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_12__5_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_12_4 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_12__4_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_11__4_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_11__5_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_12__4_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_12__4_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_12_3 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_12__3_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_11__3_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_11__4_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_12__3_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_12__3_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_12_2 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_12__2_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_11__2_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_11__3_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_12__2_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_12__2_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S2_12_1 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_12__1_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_11__1_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_11__2_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_12__1_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_12__1_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S1_12_0 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_12__0_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_11__0_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_11__1_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_12__0_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_A1_10_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S14_13 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_n86), .B(
        my_filter_adder_mult_3_multiplication_mult_21_n100), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_ab_13__13_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_13__13_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_13__13_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S5_12 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_13__12_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_12__12_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_ab_12__13_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_13__12_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_13__12_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S4_11 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_13__11_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_12__11_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_12__12_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_13__11_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_13__11_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S4_10 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_13__10_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_12__10_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_12__11_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_13__10_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_13__10_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S4_9 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_13__9_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_12__9_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_12__10_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_13__9_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_13__9_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S4_8 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_13__8_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_12__8_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_12__9_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_13__8_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_13__8_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S4_7 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_13__7_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_12__7_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_12__8_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_13__7_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_13__7_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S4_6 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_13__6_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_12__6_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_12__7_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_13__6_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_13__6_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S4_5 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_13__5_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_12__5_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_12__6_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_13__5_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_13__5_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S4_4 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_13__4_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_12__4_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_12__5_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_13__4_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_13__4_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S4_3 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_13__3_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_12__3_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_12__4_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_13__3_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_13__3_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S4_2 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_13__2_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_12__2_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_12__3_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_13__2_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_13__2_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S4_1 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_13__1_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_12__1_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_12__2_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_13__1_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_13__1_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S4_0 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_ab_13__0_), .B(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_12__0_), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_12__1_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_CARRYB_13__0_), .S(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_13__0_) );
  FA_X1 my_filter_adder_mult_3_multiplication_mult_21_S14_13_0 ( .A(
        my_filter_q_reg_chain_4__13_), .B(my_filter_q_reg_coeff[97]), .CI(
        my_filter_adder_mult_3_multiplication_mult_21_SUMB_13__0_), .CO(
        my_filter_adder_mult_3_multiplication_mult_21_A2_12_), .S(
        my_filter_adder_mult_3_res_mult[0]) );
  OAI21_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U72 ( .B1(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n15), .B2(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n16), .A(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n17), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n13) );
  NAND2_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U71 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_A2_12_), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n29), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n56) );
  OAI21_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U70 ( .B1(
        my_filter_adder_mult_3_multiplication_mult_21_A2_12_), .B2(
        my_filter_adder_mult_3_multiplication_mult_21_n29), .A(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n56), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n59) );
  INV_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U69 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n59), .ZN(
        my_filter_adder_mult_3_res_mult[1]) );
  AND2_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U68 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n51), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n48), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n20) );
  AND2_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U66 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n50), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n40), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n28) );
  AND2_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U65 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n49), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n38), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n36) );
  AND2_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U64 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n42), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n36), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n44) );
  NAND2_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U63 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n44), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n41), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n17) );
  NAND2_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U61 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n43), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n39), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n25) );
  NAND2_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U60 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n47), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n37), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n33) );
  NAND2_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U59 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n46), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n45), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n41) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U58 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n44), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n41), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n15) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U56 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n43), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n39), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n23) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U55 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n47), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n37), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n31) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U54 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n46), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n45), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n39) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U53 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n51), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n48), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n21) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U51 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n50), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n40), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n29) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U50 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n49), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n38), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n37) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U49 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n42), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n36), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n45) );
  AND2_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U48 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n35), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n30), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n52) );
  NAND2_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U46 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n34), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n32), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n49) );
  NAND2_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U45 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n33), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n31), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n57) );
  INV_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U44 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n55), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n60) );
  NAND2_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U43 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n60), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n57), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n58) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U41 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n34), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n32), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n47) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U40 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n33), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n31), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n55) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U39 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_n35), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_n30), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n53) );
  OAI21_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U38 ( .B1(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n55), .B2(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n56), .A(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n57), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n51) );
  OAI21_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U36 ( .B1(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n23), .B2(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n24), .A(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n25), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n19) );
  OAI21_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U35 ( .B1(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n31), .B2(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n32), .A(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n33), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n27) );
  INV_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U34 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n21), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n63) );
  AOI21_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U33 ( .B1(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n63), .B2(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n19), .A(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n20), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n16) );
  INV_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U31 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n29), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n71) );
  AOI21_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U30 ( .B1(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n71), .B2(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n27), .A(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n28), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n24) );
  INV_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U29 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n15), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n62) );
  NAND2_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U28 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n62), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n17), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n18) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U26 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n20), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n21), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n22) );
  INV_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U25 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n23), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n64) );
  NAND2_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U24 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n64), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n25), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n26) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U23 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n28), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n29), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n30) );
  INV_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U21 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n31), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n70) );
  NAND2_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U20 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n70), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n33), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n34) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U19 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n36), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n37), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n38) );
  INV_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U18 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n39), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n68) );
  NAND2_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U16 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n68), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n41), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n42) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U13 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n44), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n45), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n46) );
  INV_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U12 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n47), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n66) );
  NAND2_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U11 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n66), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n49), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n50) );
  NOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U10 ( .A1(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n52), .A2(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n53), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n54) );
  OAI21_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U9 ( .B1(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n39), .B2(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n40), .A(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n41), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n35) );
  OAI21_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U8 ( .B1(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n47), .B2(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n48), .A(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n49), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n43) );
  INV_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U7 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n37), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n69) );
  AOI21_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U6 ( .B1(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n69), .B2(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n35), .A(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n36), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n32) );
  INV_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U5 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n45), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n67) );
  AOI21_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U4 ( .B1(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n67), .B2(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n43), .A(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n44), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n40) );
  INV_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U3 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n53), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n65) );
  AOI21_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U2 ( .B1(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n65), .B2(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n51), .A(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n52), .ZN(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n48) );
  XOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U67 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n56), .B(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n58), .Z(
        my_filter_adder_mult_3_res_mult[2]) );
  XOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U62 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n51), .B(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n54), .Z(
        my_filter_adder_mult_3_res_mult[3]) );
  XOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U57 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n50), .B(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n48), .Z(
        my_filter_adder_mult_3_res_mult[4]) );
  XOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U52 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n43), .B(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n46), .Z(
        my_filter_adder_mult_3_res_mult[5]) );
  XOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U47 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n42), .B(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n40), .Z(
        my_filter_adder_mult_3_res_mult[6]) );
  XOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U42 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n35), .B(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n38), .Z(
        my_filter_adder_mult_3_res_mult[7]) );
  XOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U37 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n34), .B(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n32), .Z(
        my_filter_adder_mult_3_res_mult[8]) );
  XOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U32 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n27), .B(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n30), .Z(
        my_filter_adder_mult_3_res_mult[9]) );
  XOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U27 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n26), .B(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n24), .Z(
        my_filter_adder_mult_3_res_mult[10]) );
  XOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U22 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n19), .B(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n22), .Z(
        my_filter_adder_mult_3_res_mult[11]) );
  XOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U17 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n18), .B(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n16), .Z(
        my_filter_adder_mult_3_res_mult[12]) );
  XOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U15 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_n52), .B(
        my_filter_adder_mult_3_multiplication_mult_21_n27), .Z(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n14) );
  XOR2_X1 my_filter_adder_mult_3_multiplication_mult_21_FS_1_U14 ( .A(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n13), .B(
        my_filter_adder_mult_3_multiplication_mult_21_FS_1_n14), .Z(
        my_filter_adder_mult_3_res_mult[13]) );
  AND2_X1 my_filter_adder_mult_3_addition_add_19_U1 ( .A1(
        my_filter_data_sum[98]), .A2(my_filter_adder_mult_3_res_mult[0]), .ZN(
        my_filter_adder_mult_3_addition_add_19_n1) );
  XOR2_X1 my_filter_adder_mult_3_addition_add_19_U2 ( .A(
        my_filter_data_sum[98]), .B(my_filter_adder_mult_3_res_mult[0]), .Z(
        my_filter_data_sum[84]) );
  FA_X1 my_filter_adder_mult_3_addition_add_19_U1_1 ( .A(
        my_filter_adder_mult_3_res_mult[1]), .B(my_filter_data_sum[99]), .CI(
        my_filter_adder_mult_3_addition_add_19_n1), .CO(
        my_filter_adder_mult_3_addition_add_19_carry[2]), .S(
        my_filter_data_sum[85]) );
  FA_X1 my_filter_adder_mult_3_addition_add_19_U1_2 ( .A(
        my_filter_adder_mult_3_res_mult[2]), .B(my_filter_data_sum[100]), .CI(
        my_filter_adder_mult_3_addition_add_19_carry[2]), .CO(
        my_filter_adder_mult_3_addition_add_19_carry[3]), .S(
        my_filter_data_sum[86]) );
  FA_X1 my_filter_adder_mult_3_addition_add_19_U1_3 ( .A(
        my_filter_adder_mult_3_res_mult[3]), .B(my_filter_data_sum[101]), .CI(
        my_filter_adder_mult_3_addition_add_19_carry[3]), .CO(
        my_filter_adder_mult_3_addition_add_19_carry[4]), .S(
        my_filter_data_sum[87]) );
  FA_X1 my_filter_adder_mult_3_addition_add_19_U1_4 ( .A(
        my_filter_adder_mult_3_res_mult[4]), .B(my_filter_data_sum[102]), .CI(
        my_filter_adder_mult_3_addition_add_19_carry[4]), .CO(
        my_filter_adder_mult_3_addition_add_19_carry[5]), .S(
        my_filter_data_sum[88]) );
  FA_X1 my_filter_adder_mult_3_addition_add_19_U1_5 ( .A(
        my_filter_adder_mult_3_res_mult[5]), .B(my_filter_data_sum[103]), .CI(
        my_filter_adder_mult_3_addition_add_19_carry[5]), .CO(
        my_filter_adder_mult_3_addition_add_19_carry[6]), .S(
        my_filter_data_sum[89]) );
  FA_X1 my_filter_adder_mult_3_addition_add_19_U1_6 ( .A(
        my_filter_adder_mult_3_res_mult[6]), .B(my_filter_data_sum[104]), .CI(
        my_filter_adder_mult_3_addition_add_19_carry[6]), .CO(
        my_filter_adder_mult_3_addition_add_19_carry[7]), .S(
        my_filter_data_sum[90]) );
  FA_X1 my_filter_adder_mult_3_addition_add_19_U1_7 ( .A(
        my_filter_adder_mult_3_res_mult[7]), .B(my_filter_data_sum[105]), .CI(
        my_filter_adder_mult_3_addition_add_19_carry[7]), .CO(
        my_filter_adder_mult_3_addition_add_19_carry[8]), .S(
        my_filter_data_sum[91]) );
  FA_X1 my_filter_adder_mult_3_addition_add_19_U1_8 ( .A(
        my_filter_adder_mult_3_res_mult[8]), .B(my_filter_data_sum[106]), .CI(
        my_filter_adder_mult_3_addition_add_19_carry[8]), .CO(
        my_filter_adder_mult_3_addition_add_19_carry[9]), .S(
        my_filter_data_sum[92]) );
  FA_X1 my_filter_adder_mult_3_addition_add_19_U1_9 ( .A(
        my_filter_adder_mult_3_res_mult[9]), .B(my_filter_data_sum[107]), .CI(
        my_filter_adder_mult_3_addition_add_19_carry[9]), .CO(
        my_filter_adder_mult_3_addition_add_19_carry[10]), .S(
        my_filter_data_sum[93]) );
  FA_X1 my_filter_adder_mult_3_addition_add_19_U1_10 ( .A(
        my_filter_adder_mult_3_res_mult[10]), .B(my_filter_data_sum[108]), 
        .CI(my_filter_adder_mult_3_addition_add_19_carry[10]), .CO(
        my_filter_adder_mult_3_addition_add_19_carry[11]), .S(
        my_filter_data_sum[94]) );
  FA_X1 my_filter_adder_mult_3_addition_add_19_U1_11 ( .A(
        my_filter_adder_mult_3_res_mult[11]), .B(my_filter_data_sum[109]), 
        .CI(my_filter_adder_mult_3_addition_add_19_carry[11]), .CO(
        my_filter_adder_mult_3_addition_add_19_carry[12]), .S(
        my_filter_data_sum[95]) );
  FA_X1 my_filter_adder_mult_3_addition_add_19_U1_12 ( .A(
        my_filter_adder_mult_3_res_mult[12]), .B(my_filter_data_sum[110]), 
        .CI(my_filter_adder_mult_3_addition_add_19_carry[12]), .CO(
        my_filter_adder_mult_3_addition_add_19_carry[13]), .S(
        my_filter_data_sum[96]) );
  FA_X1 my_filter_adder_mult_3_addition_add_19_U1_13 ( .A(
        my_filter_adder_mult_3_res_mult[13]), .B(my_filter_data_sum[111]), 
        .CI(my_filter_adder_mult_3_addition_add_19_carry[13]), .S(
        my_filter_data_sum[97]) );
  INV_X1 my_filter_adder_mult_4_multiplication_mult_21_U276 ( .A(
        my_filter_q_reg_chain_5__12_), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_n87) );
  INV_X1 my_filter_adder_mult_4_multiplication_mult_21_U275 ( .A(
        my_filter_q_reg_chain_5__13_), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_n86) );
  AND3_X1 my_filter_adder_mult_4_multiplication_mult_21_U274 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_ab_1__1_), .A2(
        my_filter_q_reg_coeff[70]), .A3(my_filter_q_reg_chain_5__0_), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_1__0_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U273 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_12__12_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U272 ( .A1(
        my_filter_q_reg_chain_5__11_), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_11__13_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U271 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_11__12_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U270 ( .A1(
        my_filter_q_reg_chain_5__10_), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_10__13_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U269 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_10__12_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U268 ( .A1(
        my_filter_q_reg_chain_5__9_), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_9__13_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U267 ( .A1(
        my_filter_q_reg_chain_5__8_), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_8__13_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U266 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n101), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_9__12_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U265 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_8__12_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U264 ( .A1(
        my_filter_q_reg_chain_5__7_), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_7__13_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U263 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_7__12_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U262 ( .A1(
        my_filter_q_reg_chain_5__6_), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_6__13_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U261 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_6__12_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U260 ( .A1(
        my_filter_q_reg_chain_5__5_), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_5__13_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U259 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_5__12_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U258 ( .A1(
        my_filter_q_reg_chain_5__4_), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_4__13_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U257 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_4__12_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U256 ( .A1(
        my_filter_q_reg_chain_5__3_), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_3__13_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U255 ( .A1(
        my_filter_q_reg_coeff[80]), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_13__10_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U254 ( .A1(
        my_filter_q_reg_coeff[81]), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_13__11_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U253 ( .A1(
        my_filter_q_reg_coeff[78]), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_13__8_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U252 ( .A1(
        my_filter_q_reg_coeff[79]), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_13__9_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U251 ( .A1(
        my_filter_q_reg_coeff[76]), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_13__6_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U250 ( .A1(
        my_filter_q_reg_coeff[77]), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_13__7_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U249 ( .A1(
        my_filter_q_reg_coeff[74]), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_13__4_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U248 ( .A1(
        my_filter_q_reg_coeff[75]), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_13__5_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U247 ( .A1(
        my_filter_q_reg_coeff[73]), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_13__3_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U246 ( .A1(
        my_filter_q_reg_coeff[82]), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_13__12_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U245 ( .A1(
        my_filter_q_reg_chain_5__12_), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_12__13_) );
  INV_X1 my_filter_adder_mult_4_multiplication_mult_21_U244 ( .A(
        my_filter_q_reg_coeff[70]), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_n113) );
  INV_X1 my_filter_adder_mult_4_multiplication_mult_21_U243 ( .A(
        my_filter_q_reg_coeff[71]), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_n112) );
  INV_X1 my_filter_adder_mult_4_multiplication_mult_21_U242 ( .A(
        my_filter_q_reg_chain_5__9_), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_n90) );
  INV_X1 my_filter_adder_mult_4_multiplication_mult_21_U241 ( .A(
        my_filter_q_reg_coeff[72]), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_n111) );
  INV_X1 my_filter_adder_mult_4_multiplication_mult_21_U240 ( .A(
        my_filter_q_reg_chain_5__11_), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_n88) );
  INV_X1 my_filter_adder_mult_4_multiplication_mult_21_U239 ( .A(
        my_filter_q_reg_chain_5__10_), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_n89) );
  INV_X1 my_filter_adder_mult_4_multiplication_mult_21_U238 ( .A(
        my_filter_q_reg_chain_5__8_), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_n91) );
  INV_X1 my_filter_adder_mult_4_multiplication_mult_21_U237 ( .A(
        my_filter_q_reg_chain_5__7_), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_n92) );
  INV_X1 my_filter_adder_mult_4_multiplication_mult_21_U236 ( .A(
        my_filter_q_reg_chain_5__6_), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_n93) );
  INV_X1 my_filter_adder_mult_4_multiplication_mult_21_U235 ( .A(
        my_filter_q_reg_chain_5__5_), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_n94) );
  INV_X1 my_filter_adder_mult_4_multiplication_mult_21_U234 ( .A(
        my_filter_q_reg_chain_5__4_), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_n95) );
  AND2_X1 my_filter_adder_mult_4_multiplication_mult_21_U233 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_ab_0__13_), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_ab_1__12_), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_n15) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U232 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_2__12_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U231 ( .A1(
        my_filter_q_reg_chain_5__1_), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_1__13_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U230 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_12__0_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U229 ( .A1(
        my_filter_q_reg_coeff[70]), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_13__0_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U228 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_3__12_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U227 ( .A1(
        my_filter_q_reg_chain_5__2_), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_2__13_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U226 ( .A1(
        my_filter_q_reg_coeff[71]), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_13__1_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U225 ( .A1(
        my_filter_q_reg_coeff[72]), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_13__2_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U224 ( .A1(
        my_filter_q_reg_chain_5__0_), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_0__13_) );
  INV_X1 my_filter_adder_mult_4_multiplication_mult_21_U223 ( .A(
        my_filter_q_reg_coeff[83]), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_n100) );
  INV_X1 my_filter_adder_mult_4_multiplication_mult_21_U222 ( .A(
        my_filter_q_reg_chain_5__0_), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_n99) );
  INV_X1 my_filter_adder_mult_4_multiplication_mult_21_U221 ( .A(
        my_filter_q_reg_chain_5__1_), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_n98) );
  INV_X1 my_filter_adder_mult_4_multiplication_mult_21_U220 ( .A(
        my_filter_q_reg_coeff[82]), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_n101) );
  INV_X1 my_filter_adder_mult_4_multiplication_mult_21_U219 ( .A(
        my_filter_q_reg_coeff[80]), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_n103) );
  INV_X1 my_filter_adder_mult_4_multiplication_mult_21_U218 ( .A(
        my_filter_q_reg_coeff[81]), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_n102) );
  INV_X1 my_filter_adder_mult_4_multiplication_mult_21_U217 ( .A(
        my_filter_q_reg_coeff[78]), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_n105) );
  INV_X1 my_filter_adder_mult_4_multiplication_mult_21_U216 ( .A(
        my_filter_q_reg_coeff[79]), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_n104) );
  INV_X1 my_filter_adder_mult_4_multiplication_mult_21_U215 ( .A(
        my_filter_q_reg_coeff[75]), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_n108) );
  INV_X1 my_filter_adder_mult_4_multiplication_mult_21_U214 ( .A(
        my_filter_q_reg_coeff[76]), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_n107) );
  INV_X1 my_filter_adder_mult_4_multiplication_mult_21_U213 ( .A(
        my_filter_q_reg_coeff[77]), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_n106) );
  INV_X1 my_filter_adder_mult_4_multiplication_mult_21_U212 ( .A(
        my_filter_q_reg_coeff[73]), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_n110) );
  INV_X1 my_filter_adder_mult_4_multiplication_mult_21_U211 ( .A(
        my_filter_q_reg_coeff[74]), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_n109) );
  INV_X1 my_filter_adder_mult_4_multiplication_mult_21_U210 ( .A(
        my_filter_q_reg_chain_5__2_), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_n97) );
  INV_X1 my_filter_adder_mult_4_multiplication_mult_21_U209 ( .A(
        my_filter_q_reg_chain_5__3_), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_n96) );
  AND2_X1 my_filter_adder_mult_4_multiplication_mult_21_U208 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_13__12_), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_13__13_), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_n3) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U207 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n100), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_13__13_) );
  AND2_X1 my_filter_adder_mult_4_multiplication_mult_21_U206 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_13__11_), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_13__12_), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_n52) );
  AND2_X1 my_filter_adder_mult_4_multiplication_mult_21_U205 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_13__9_), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_13__10_), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_n50) );
  AND2_X1 my_filter_adder_mult_4_multiplication_mult_21_U204 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_13__7_), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_13__8_), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_n49) );
  AND2_X1 my_filter_adder_mult_4_multiplication_mult_21_U203 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_13__5_), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_13__6_), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_n48) );
  AND2_X1 my_filter_adder_mult_4_multiplication_mult_21_U202 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_13__3_), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_13__4_), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_n40) );
  AND2_X1 my_filter_adder_mult_4_multiplication_mult_21_U201 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_13__1_), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_13__2_), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_n32) );
  AND2_X1 my_filter_adder_mult_4_multiplication_mult_21_U200 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_13__10_), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_13__11_), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_n43) );
  AND2_X1 my_filter_adder_mult_4_multiplication_mult_21_U199 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_13__8_), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_13__9_), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_n42) );
  AND2_X1 my_filter_adder_mult_4_multiplication_mult_21_U198 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_13__6_), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_13__7_), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_n41) );
  AND2_X1 my_filter_adder_mult_4_multiplication_mult_21_U197 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_13__4_), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_13__5_), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_n39) );
  AND2_X1 my_filter_adder_mult_4_multiplication_mult_21_U196 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_13__2_), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_13__3_), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_n46) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U195 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_12__11_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U194 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_12__9_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U193 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_12__10_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U192 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_11__10_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U191 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_11__11_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U190 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_12__7_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U189 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_12__8_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U188 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_10__11_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U187 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_11__8_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U186 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_11__9_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U185 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_12__5_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U184 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_12__6_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U183 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_10__9_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U182 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_10__10_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U181 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_11__6_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U180 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_11__7_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U179 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n103), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_9__10_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U178 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n102), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_9__11_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U177 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_12__4_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U176 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_10__7_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U175 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_10__8_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U174 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_8__11_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U173 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_11__5_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U172 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n105), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_9__8_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U171 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n104), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_9__9_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U170 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_10__6_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U169 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_8__9_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U168 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_8__10_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U167 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n106), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_9__7_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U166 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_7__10_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U165 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_7__11_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U164 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_8__8_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U163 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_6__11_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U162 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_7__9_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U161 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_6__10_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U160 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_5__11_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U159 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_0__2_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U158 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n98), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n112), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_1__1_) );
  AND2_X1 my_filter_adder_mult_4_multiplication_mult_21_U157 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_13__0_), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_13__1_), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_n31) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U156 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_12__1_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U155 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_10__0_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U154 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_11__0_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U153 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_11__1_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U152 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_10__1_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U151 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_8__0_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U150 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n113), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_9__0_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U149 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n112), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_9__1_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U148 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n110), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_9__3_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U147 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_8__1_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U146 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_8__3_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U145 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_6__0_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U144 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_7__0_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U143 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_7__1_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U142 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_7__3_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U141 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_7__4_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U140 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_7__5_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U139 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_6__1_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U138 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_6__3_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U137 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_6__5_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U136 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_4__0_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U135 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_5__0_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U134 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_5__1_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U133 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_5__3_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U132 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_5__4_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U131 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_5__5_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U130 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_5__6_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U129 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_5__7_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U128 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_4__1_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U127 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_4__3_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U126 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_4__5_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U125 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_2__0_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U124 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_3__0_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U123 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_3__1_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U122 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_3__3_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U121 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_3__4_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U120 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_3__5_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U119 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_3__6_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U118 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_3__7_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U117 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_3__8_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U116 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_3__9_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U115 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_12__2_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U114 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_12__3_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U113 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_11__3_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U112 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_11__4_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U111 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_10__4_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U110 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_10__5_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U109 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_11__2_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U108 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n108), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_9__5_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U107 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n107), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_9__6_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U106 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_10__2_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U105 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_10__3_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U104 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_8__6_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U103 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_8__7_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U102 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n111), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_9__2_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U101 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n109), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_9__4_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U100 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_7__7_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U99 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_7__8_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U98 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_8__2_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U97 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_8__4_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U96 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_8__5_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U95 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_6__8_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U94 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_6__9_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U93 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_7__2_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U92 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_7__6_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U91 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_5__9_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U90 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_5__10_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U89 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_6__2_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U88 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_6__4_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U87 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_6__6_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U86 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_6__7_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U85 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_4__10_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U84 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_4__11_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U83 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_5__2_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U82 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_5__8_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U81 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_3__11_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U80 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_4__2_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U79 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_4__4_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U78 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_4__6_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U77 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_4__7_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U76 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_4__8_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U75 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_4__9_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U74 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_3__2_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U73 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_3__10_) );
  AND2_X1 my_filter_adder_mult_4_multiplication_mult_21_U72 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_ab_0__2_), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_ab_1__1_), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_n14) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U71 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_2__1_) );
  AND2_X1 my_filter_adder_mult_4_multiplication_mult_21_U70 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_ab_0__3_), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_ab_1__2_), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_n13) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U69 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_2__2_) );
  AND2_X1 my_filter_adder_mult_4_multiplication_mult_21_U68 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_ab_0__4_), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_ab_1__3_), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_n12) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U67 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_2__3_) );
  AND2_X1 my_filter_adder_mult_4_multiplication_mult_21_U66 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_ab_0__5_), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_ab_1__4_), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_n11) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U65 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_2__4_) );
  AND2_X1 my_filter_adder_mult_4_multiplication_mult_21_U64 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_ab_0__6_), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_ab_1__5_), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_n22) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U63 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_2__5_) );
  AND2_X1 my_filter_adder_mult_4_multiplication_mult_21_U62 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_ab_0__7_), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_ab_1__6_), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_n21) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U61 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_2__6_) );
  AND2_X1 my_filter_adder_mult_4_multiplication_mult_21_U60 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_ab_0__8_), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_ab_1__7_), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_n4) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U59 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_2__7_) );
  AND2_X1 my_filter_adder_mult_4_multiplication_mult_21_U58 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_ab_0__9_), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_ab_1__8_), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_n8) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U57 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_2__8_) );
  AND2_X1 my_filter_adder_mult_4_multiplication_mult_21_U56 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_ab_0__10_), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_ab_1__9_), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_n7) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U55 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_2__9_) );
  AND2_X1 my_filter_adder_mult_4_multiplication_mult_21_U54 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_ab_0__11_), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_ab_1__10_), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_n6) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U52 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_2__10_) );
  AND2_X1 my_filter_adder_mult_4_multiplication_mult_21_U50 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_ab_0__12_), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_ab_1__11_), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_n5) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U49 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_2__11_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U48 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_1__12_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U46 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_1__2_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U43 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_1__3_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U42 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_1__4_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U41 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_1__5_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U40 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_1__6_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U39 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_1__7_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U32 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_1__8_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U31 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_1__9_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U21 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_1__10_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U20 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_1__11_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U14 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_0__3_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U13 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_0__4_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U12 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_0__5_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U11 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_0__6_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U10 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_0__7_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U7 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_0__8_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U6 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_0__9_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U5 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_0__10_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U4 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_0__11_) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U3 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_ab_0__12_) );
  INV_X1 my_filter_adder_mult_4_multiplication_mult_21_U2 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_13__13_), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_n85) );
  XOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U51 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_13__12_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_13__13_), .Z(
        my_filter_adder_mult_4_multiplication_mult_21_n51) );
  XOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U47 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_13__10_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_13__11_), .Z(
        my_filter_adder_mult_4_multiplication_mult_21_n47) );
  XOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U45 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_13__5_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_13__6_), .Z(
        my_filter_adder_mult_4_multiplication_mult_21_n45) );
  XOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U44 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_13__3_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_13__4_), .Z(
        my_filter_adder_mult_4_multiplication_mult_21_n44) );
  XOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U38 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_13__11_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_13__12_), .Z(
        my_filter_adder_mult_4_multiplication_mult_21_n38) );
  XOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U37 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_13__8_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_13__9_), .Z(
        my_filter_adder_mult_4_multiplication_mult_21_n37) );
  XOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U36 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_13__9_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_13__10_), .Z(
        my_filter_adder_mult_4_multiplication_mult_21_n36) );
  XOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U35 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_13__6_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_13__7_), .Z(
        my_filter_adder_mult_4_multiplication_mult_21_n35) );
  XOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U34 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_13__7_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_13__8_), .Z(
        my_filter_adder_mult_4_multiplication_mult_21_n34) );
  XOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U33 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_13__4_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_13__5_), .Z(
        my_filter_adder_mult_4_multiplication_mult_21_n33) );
  XOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U30 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_13__1_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_13__2_), .Z(
        my_filter_adder_mult_4_multiplication_mult_21_n30) );
  XOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U29 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_13__2_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_13__3_), .Z(
        my_filter_adder_mult_4_multiplication_mult_21_n29) );
  XOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U28 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_13__0_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_13__1_), .Z(
        my_filter_adder_mult_4_multiplication_mult_21_n28) );
  XOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U26 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_1__1_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_ab_0__2_), .Z(
        my_filter_adder_mult_4_multiplication_mult_21_n27) );
  XOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U25 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_1__2_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_ab_0__3_), .Z(
        my_filter_adder_mult_4_multiplication_mult_21_n26) );
  XOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U24 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_1__3_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_ab_0__4_), .Z(
        my_filter_adder_mult_4_multiplication_mult_21_n25) );
  XOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U23 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_1__4_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_ab_0__5_), .Z(
        my_filter_adder_mult_4_multiplication_mult_21_n24) );
  XOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U22 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_1__5_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_ab_0__6_), .Z(
        my_filter_adder_mult_4_multiplication_mult_21_n23) );
  XOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U19 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_1__12_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_ab_0__13_), .Z(
        my_filter_adder_mult_4_multiplication_mult_21_n20) );
  XOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U18 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_1__8_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_ab_0__9_), .Z(
        my_filter_adder_mult_4_multiplication_mult_21_n19) );
  XOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U17 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_1__9_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_ab_0__10_), .Z(
        my_filter_adder_mult_4_multiplication_mult_21_n18) );
  XOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U16 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_1__10_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_ab_0__11_), .Z(
        my_filter_adder_mult_4_multiplication_mult_21_n17) );
  XOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U15 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_1__11_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_ab_0__12_), .Z(
        my_filter_adder_mult_4_multiplication_mult_21_n16) );
  XOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U9 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_1__6_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_ab_0__7_), .Z(
        my_filter_adder_mult_4_multiplication_mult_21_n10) );
  XOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_U8 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_1__7_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_ab_0__8_), .Z(
        my_filter_adder_mult_4_multiplication_mult_21_n9) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S3_2_12 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_2__12_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_n15), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_ab_1__13_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_2__12_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_2__12_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_2_11 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_2__11_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_n5), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_n20), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_2__11_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_2__11_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_2_10 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_2__10_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_n6), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_n16), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_2__10_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_2__10_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_2_9 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_2__9_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_n7), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_n17), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_2__9_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_2__9_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_2_8 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_2__8_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_n8), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_n18), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_2__8_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_2__8_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_2_7 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_2__7_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_n4), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_n19), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_2__7_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_2__7_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_2_6 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_2__6_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_n21), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_n9), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_2__6_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_2__6_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_2_5 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_2__5_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_n22), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_n10), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_2__5_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_2__5_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_2_4 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_2__4_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_n11), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_n23), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_2__4_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_2__4_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_2_3 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_2__3_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_n12), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_n24), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_2__3_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_2__3_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_2_2 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_2__2_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_n13), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_n25), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_2__2_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_2__2_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_2_1 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_2__1_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_n14), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_n26), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_2__1_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_2__1_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S1_2_0 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_2__0_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_1__0_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_n27), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_2__0_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_A1_0_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S3_3_12 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_3__12_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_2__12_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_ab_2__13_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_3__12_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_3__12_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_3_11 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_3__11_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_2__11_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_2__12_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_3__11_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_3__11_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_3_10 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_3__10_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_2__10_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_2__11_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_3__10_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_3__10_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_3_9 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_3__9_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_2__9_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_2__10_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_3__9_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_3__9_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_3_8 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_3__8_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_2__8_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_2__9_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_3__8_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_3__8_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_3_7 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_3__7_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_2__7_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_2__8_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_3__7_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_3__7_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_3_6 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_3__6_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_2__6_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_2__7_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_3__6_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_3__6_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_3_5 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_3__5_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_2__5_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_2__6_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_3__5_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_3__5_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_3_4 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_3__4_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_2__4_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_2__5_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_3__4_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_3__4_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_3_3 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_3__3_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_2__3_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_2__4_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_3__3_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_3__3_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_3_2 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_3__2_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_2__2_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_2__3_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_3__2_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_3__2_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_3_1 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_3__1_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_2__1_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_2__2_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_3__1_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_3__1_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S1_3_0 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_3__0_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_2__0_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_2__1_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_3__0_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_A1_1_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S3_4_12 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_4__12_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_3__12_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_ab_3__13_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_4__12_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_4__12_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_4_11 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_4__11_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_3__11_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_3__12_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_4__11_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_4__11_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_4_10 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_4__10_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_3__10_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_3__11_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_4__10_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_4__10_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_4_9 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_4__9_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_3__9_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_3__10_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_4__9_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_4__9_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_4_8 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_4__8_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_3__8_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_3__9_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_4__8_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_4__8_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_4_7 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_4__7_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_3__7_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_3__8_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_4__7_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_4__7_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_4_6 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_4__6_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_3__6_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_3__7_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_4__6_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_4__6_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_4_5 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_4__5_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_3__5_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_3__6_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_4__5_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_4__5_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_4_4 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_4__4_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_3__4_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_3__5_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_4__4_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_4__4_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_4_3 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_4__3_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_3__3_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_3__4_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_4__3_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_4__3_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_4_2 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_4__2_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_3__2_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_3__3_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_4__2_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_4__2_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_4_1 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_4__1_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_3__1_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_3__2_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_4__1_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_4__1_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S1_4_0 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_4__0_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_3__0_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_3__1_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_4__0_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_A1_2_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S3_5_12 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_5__12_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_4__12_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_ab_4__13_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_5__12_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_5__12_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_5_11 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_5__11_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_4__11_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_4__12_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_5__11_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_5__11_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_5_10 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_5__10_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_4__10_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_4__11_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_5__10_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_5__10_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_5_9 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_5__9_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_4__9_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_4__10_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_5__9_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_5__9_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_5_8 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_5__8_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_4__8_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_4__9_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_5__8_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_5__8_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_5_7 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_5__7_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_4__7_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_4__8_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_5__7_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_5__7_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_5_6 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_5__6_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_4__6_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_4__7_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_5__6_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_5__6_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_5_5 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_5__5_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_4__5_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_4__6_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_5__5_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_5__5_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_5_4 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_5__4_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_4__4_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_4__5_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_5__4_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_5__4_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_5_3 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_5__3_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_4__3_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_4__4_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_5__3_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_5__3_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_5_2 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_5__2_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_4__2_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_4__3_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_5__2_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_5__2_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_5_1 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_5__1_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_4__1_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_4__2_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_5__1_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_5__1_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S1_5_0 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_5__0_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_4__0_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_4__1_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_5__0_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_A1_3_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S3_6_12 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_6__12_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_5__12_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_ab_5__13_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_6__12_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_6__12_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_6_11 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_6__11_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_5__11_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_5__12_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_6__11_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_6__11_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_6_10 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_6__10_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_5__10_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_5__11_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_6__10_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_6__10_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_6_9 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_6__9_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_5__9_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_5__10_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_6__9_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_6__9_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_6_8 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_6__8_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_5__8_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_5__9_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_6__8_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_6__8_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_6_7 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_6__7_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_5__7_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_5__8_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_6__7_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_6__7_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_6_6 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_6__6_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_5__6_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_5__7_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_6__6_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_6__6_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_6_5 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_6__5_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_5__5_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_5__6_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_6__5_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_6__5_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_6_4 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_6__4_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_5__4_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_5__5_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_6__4_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_6__4_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_6_3 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_6__3_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_5__3_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_5__4_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_6__3_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_6__3_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_6_2 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_6__2_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_5__2_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_5__3_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_6__2_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_6__2_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_6_1 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_6__1_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_5__1_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_5__2_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_6__1_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_6__1_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S1_6_0 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_6__0_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_5__0_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_5__1_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_6__0_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_A1_4_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S3_7_12 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_7__12_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_6__12_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_ab_6__13_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_7__12_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_7__12_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_7_11 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_7__11_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_6__11_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_6__12_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_7__11_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_7__11_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_7_10 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_7__10_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_6__10_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_6__11_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_7__10_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_7__10_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_7_9 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_7__9_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_6__9_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_6__10_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_7__9_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_7__9_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_7_8 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_7__8_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_6__8_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_6__9_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_7__8_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_7__8_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_7_7 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_7__7_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_6__7_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_6__8_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_7__7_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_7__7_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_7_6 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_7__6_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_6__6_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_6__7_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_7__6_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_7__6_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_7_5 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_7__5_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_6__5_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_6__6_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_7__5_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_7__5_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_7_4 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_7__4_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_6__4_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_6__5_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_7__4_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_7__4_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_7_3 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_7__3_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_6__3_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_6__4_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_7__3_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_7__3_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_7_2 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_7__2_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_6__2_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_6__3_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_7__2_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_7__2_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_7_1 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_7__1_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_6__1_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_6__2_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_7__1_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_7__1_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S1_7_0 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_7__0_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_6__0_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_6__1_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_7__0_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_A1_5_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S3_8_12 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_8__12_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_7__12_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_ab_7__13_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_8__12_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_8__12_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_8_11 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_8__11_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_7__11_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_7__12_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_8__11_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_8__11_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_8_10 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_8__10_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_7__10_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_7__11_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_8__10_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_8__10_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_8_9 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_8__9_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_7__9_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_7__10_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_8__9_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_8__9_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_8_8 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_8__8_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_7__8_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_7__9_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_8__8_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_8__8_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_8_7 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_8__7_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_7__7_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_7__8_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_8__7_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_8__7_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_8_6 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_8__6_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_7__6_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_7__7_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_8__6_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_8__6_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_8_5 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_8__5_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_7__5_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_7__6_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_8__5_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_8__5_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_8_4 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_8__4_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_7__4_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_7__5_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_8__4_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_8__4_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_8_3 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_8__3_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_7__3_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_7__4_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_8__3_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_8__3_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_8_2 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_8__2_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_7__2_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_7__3_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_8__2_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_8__2_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_8_1 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_8__1_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_7__1_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_7__2_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_8__1_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_8__1_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S1_8_0 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_8__0_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_7__0_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_7__1_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_8__0_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_A1_6_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S3_9_12 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_9__12_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_8__12_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_ab_8__13_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_9__12_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_9__12_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_9_11 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_9__11_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_8__11_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_8__12_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_9__11_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_9__11_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_9_10 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_9__10_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_8__10_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_8__11_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_9__10_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_9__10_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_9_9 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_9__9_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_8__9_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_8__10_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_9__9_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_9__9_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_9_8 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_9__8_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_8__8_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_8__9_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_9__8_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_9__8_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_9_7 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_9__7_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_8__7_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_8__8_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_9__7_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_9__7_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_9_6 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_9__6_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_8__6_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_8__7_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_9__6_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_9__6_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_9_5 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_9__5_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_8__5_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_8__6_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_9__5_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_9__5_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_9_4 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_9__4_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_8__4_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_8__5_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_9__4_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_9__4_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_9_3 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_9__3_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_8__3_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_8__4_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_9__3_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_9__3_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_9_2 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_9__2_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_8__2_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_8__3_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_9__2_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_9__2_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_9_1 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_9__1_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_8__1_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_8__2_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_9__1_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_9__1_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S1_9_0 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_9__0_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_8__0_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_8__1_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_9__0_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_A1_7_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S3_10_12 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_10__12_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_9__12_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_ab_9__13_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_10__12_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_10__12_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_10_11 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_10__11_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_9__11_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_9__12_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_10__11_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_10__11_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_10_10 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_10__10_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_9__10_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_9__11_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_10__10_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_10__10_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_10_9 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_10__9_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_9__9_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_9__10_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_10__9_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_10__9_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_10_8 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_10__8_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_9__8_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_9__9_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_10__8_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_10__8_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_10_7 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_10__7_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_9__7_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_9__8_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_10__7_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_10__7_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_10_6 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_10__6_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_9__6_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_9__7_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_10__6_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_10__6_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_10_5 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_10__5_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_9__5_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_9__6_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_10__5_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_10__5_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_10_4 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_10__4_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_9__4_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_9__5_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_10__4_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_10__4_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_10_3 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_10__3_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_9__3_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_9__4_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_10__3_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_10__3_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_10_2 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_10__2_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_9__2_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_9__3_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_10__2_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_10__2_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_10_1 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_10__1_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_9__1_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_9__2_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_10__1_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_10__1_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S1_10_0 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_10__0_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_9__0_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_9__1_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_10__0_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_A1_8_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S3_11_12 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_11__12_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_10__12_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_ab_10__13_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_11__12_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_11__12_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_11_11 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_11__11_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_10__11_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_10__12_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_11__11_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_11__11_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_11_10 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_11__10_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_10__10_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_10__11_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_11__10_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_11__10_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_11_9 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_11__9_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_10__9_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_10__10_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_11__9_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_11__9_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_11_8 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_11__8_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_10__8_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_10__9_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_11__8_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_11__8_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_11_7 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_11__7_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_10__7_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_10__8_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_11__7_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_11__7_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_11_6 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_11__6_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_10__6_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_10__7_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_11__6_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_11__6_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_11_5 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_11__5_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_10__5_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_10__6_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_11__5_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_11__5_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_11_4 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_11__4_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_10__4_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_10__5_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_11__4_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_11__4_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_11_3 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_11__3_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_10__3_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_10__4_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_11__3_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_11__3_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_11_2 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_11__2_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_10__2_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_10__3_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_11__2_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_11__2_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_11_1 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_11__1_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_10__1_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_10__2_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_11__1_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_11__1_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S1_11_0 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_11__0_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_10__0_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_10__1_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_11__0_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_A1_9_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S3_12_12 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_12__12_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_11__12_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_ab_11__13_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_12__12_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_12__12_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_12_11 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_12__11_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_11__11_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_11__12_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_12__11_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_12__11_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_12_10 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_12__10_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_11__10_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_11__11_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_12__10_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_12__10_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_12_9 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_12__9_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_11__9_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_11__10_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_12__9_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_12__9_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_12_8 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_12__8_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_11__8_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_11__9_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_12__8_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_12__8_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_12_7 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_12__7_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_11__7_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_11__8_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_12__7_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_12__7_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_12_6 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_12__6_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_11__6_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_11__7_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_12__6_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_12__6_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_12_5 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_12__5_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_11__5_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_11__6_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_12__5_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_12__5_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_12_4 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_12__4_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_11__4_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_11__5_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_12__4_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_12__4_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_12_3 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_12__3_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_11__3_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_11__4_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_12__3_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_12__3_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_12_2 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_12__2_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_11__2_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_11__3_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_12__2_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_12__2_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S2_12_1 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_12__1_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_11__1_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_11__2_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_12__1_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_12__1_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S1_12_0 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_12__0_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_11__0_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_11__1_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_12__0_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_A1_10_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S14_13 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_n86), .B(
        my_filter_adder_mult_4_multiplication_mult_21_n100), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_ab_13__13_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_13__13_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_13__13_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S5_12 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_13__12_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_12__12_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_ab_12__13_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_13__12_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_13__12_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S4_11 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_13__11_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_12__11_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_12__12_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_13__11_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_13__11_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S4_10 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_13__10_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_12__10_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_12__11_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_13__10_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_13__10_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S4_9 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_13__9_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_12__9_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_12__10_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_13__9_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_13__9_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S4_8 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_13__8_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_12__8_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_12__9_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_13__8_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_13__8_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S4_7 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_13__7_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_12__7_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_12__8_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_13__7_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_13__7_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S4_6 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_13__6_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_12__6_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_12__7_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_13__6_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_13__6_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S4_5 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_13__5_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_12__5_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_12__6_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_13__5_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_13__5_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S4_4 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_13__4_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_12__4_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_12__5_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_13__4_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_13__4_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S4_3 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_13__3_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_12__3_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_12__4_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_13__3_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_13__3_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S4_2 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_13__2_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_12__2_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_12__3_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_13__2_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_13__2_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S4_1 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_13__1_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_12__1_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_12__2_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_13__1_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_13__1_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S4_0 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_ab_13__0_), .B(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_12__0_), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_12__1_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_CARRYB_13__0_), .S(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_13__0_) );
  FA_X1 my_filter_adder_mult_4_multiplication_mult_21_S14_13_0 ( .A(
        my_filter_q_reg_chain_5__13_), .B(my_filter_q_reg_coeff[83]), .CI(
        my_filter_adder_mult_4_multiplication_mult_21_SUMB_13__0_), .CO(
        my_filter_adder_mult_4_multiplication_mult_21_A2_12_), .S(
        my_filter_adder_mult_4_res_mult[0]) );
  NAND2_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U72 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_A2_12_), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n28), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n56) );
  OAI21_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U71 ( .B1(
        my_filter_adder_mult_4_multiplication_mult_21_A2_12_), .B2(
        my_filter_adder_mult_4_multiplication_mult_21_n28), .A(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n56), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n59) );
  INV_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U70 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n59), .ZN(
        my_filter_adder_mult_4_res_mult[1]) );
  AND2_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U69 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n50), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n47), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n20) );
  AND2_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U68 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n49), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n37), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n28) );
  AND2_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U66 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n48), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n35), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n36) );
  AND2_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U65 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n40), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n33), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n44) );
  AND2_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U64 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n32), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n29), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n52) );
  NAND2_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U63 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n43), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n38), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n17) );
  NAND2_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U61 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n42), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n36), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n25) );
  NAND2_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U60 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n41), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n34), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n33) );
  NAND2_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U59 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n39), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n45), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n41) );
  NAND2_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U58 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n46), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n44), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n49) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U56 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n43), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n38), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n15) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U55 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n42), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n36), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n23) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U54 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n41), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n34), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n31) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U53 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n39), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n45), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n39) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U51 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n46), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n44), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n47) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U50 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n50), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n47), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n21) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U49 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n49), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n37), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n29) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U48 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n48), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n35), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n37) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U46 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n40), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n33), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n45) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U45 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n32), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n29), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n53) );
  NAND2_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U44 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n31), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n30), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n57) );
  INV_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U43 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n55), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n60) );
  NAND2_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U41 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n60), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n57), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n58) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U40 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_n31), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_n30), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n55) );
  OAI21_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U39 ( .B1(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n55), .B2(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n56), .A(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n57), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n51) );
  OAI21_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U38 ( .B1(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n15), .B2(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n16), .A(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n17), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n13) );
  OAI21_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U36 ( .B1(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n23), .B2(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n24), .A(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n25), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n19) );
  OAI21_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U35 ( .B1(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n31), .B2(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n32), .A(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n33), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n27) );
  OAI21_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U34 ( .B1(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n39), .B2(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n40), .A(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n41), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n35) );
  OAI21_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U33 ( .B1(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n47), .B2(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n48), .A(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n49), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n43) );
  INV_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U31 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n21), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n63) );
  AOI21_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U30 ( .B1(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n63), .B2(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n19), .A(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n20), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n16) );
  INV_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U29 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n29), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n71) );
  AOI21_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U28 ( .B1(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n71), .B2(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n27), .A(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n28), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n24) );
  INV_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U26 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n37), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n69) );
  AOI21_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U25 ( .B1(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n69), .B2(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n35), .A(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n36), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n32) );
  INV_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U24 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n45), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n67) );
  AOI21_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U23 ( .B1(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n67), .B2(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n43), .A(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n44), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n40) );
  INV_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U21 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n15), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n62) );
  NAND2_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U20 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n62), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n17), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n18) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U19 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n20), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n21), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n22) );
  INV_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U18 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n23), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n64) );
  NAND2_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U16 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n64), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n25), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n26) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U13 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n28), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n29), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n30) );
  INV_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U12 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n31), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n70) );
  NAND2_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U11 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n70), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n33), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n34) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U10 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n36), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n37), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n38) );
  INV_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U9 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n39), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n68) );
  NAND2_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U8 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n68), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n41), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n42) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U7 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n44), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n45), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n46) );
  INV_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U6 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n47), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n66) );
  NAND2_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U5 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n66), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n49), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n50) );
  NOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U4 ( .A1(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n52), .A2(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n53), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n54) );
  INV_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U3 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n53), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n65) );
  AOI21_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U2 ( .B1(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n65), .B2(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n51), .A(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n52), .ZN(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n48) );
  XOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U67 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n56), .B(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n58), .Z(
        my_filter_adder_mult_4_res_mult[2]) );
  XOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U62 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n51), .B(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n54), .Z(
        my_filter_adder_mult_4_res_mult[3]) );
  XOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U57 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n50), .B(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n48), .Z(
        my_filter_adder_mult_4_res_mult[4]) );
  XOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U52 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n43), .B(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n46), .Z(
        my_filter_adder_mult_4_res_mult[5]) );
  XOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U47 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n42), .B(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n40), .Z(
        my_filter_adder_mult_4_res_mult[6]) );
  XOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U42 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n35), .B(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n38), .Z(
        my_filter_adder_mult_4_res_mult[7]) );
  XOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U37 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n34), .B(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n32), .Z(
        my_filter_adder_mult_4_res_mult[8]) );
  XOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U32 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n27), .B(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n30), .Z(
        my_filter_adder_mult_4_res_mult[9]) );
  XOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U27 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n26), .B(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n24), .Z(
        my_filter_adder_mult_4_res_mult[10]) );
  XOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U22 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n19), .B(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n22), .Z(
        my_filter_adder_mult_4_res_mult[11]) );
  XOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U17 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n18), .B(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n16), .Z(
        my_filter_adder_mult_4_res_mult[12]) );
  XOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U15 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_n52), .B(
        my_filter_adder_mult_4_multiplication_mult_21_n51), .Z(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n14) );
  XOR2_X1 my_filter_adder_mult_4_multiplication_mult_21_FS_1_U14 ( .A(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n13), .B(
        my_filter_adder_mult_4_multiplication_mult_21_FS_1_n14), .Z(
        my_filter_adder_mult_4_res_mult[13]) );
  AND2_X1 my_filter_adder_mult_4_addition_add_19_U1 ( .A1(
        my_filter_data_sum[84]), .A2(my_filter_adder_mult_4_res_mult[0]), .ZN(
        my_filter_adder_mult_4_addition_add_19_n1) );
  XOR2_X1 my_filter_adder_mult_4_addition_add_19_U2 ( .A(
        my_filter_data_sum[84]), .B(my_filter_adder_mult_4_res_mult[0]), .Z(
        my_filter_data_sum[70]) );
  FA_X1 my_filter_adder_mult_4_addition_add_19_U1_1 ( .A(
        my_filter_adder_mult_4_res_mult[1]), .B(my_filter_data_sum[85]), .CI(
        my_filter_adder_mult_4_addition_add_19_n1), .CO(
        my_filter_adder_mult_4_addition_add_19_carry[2]), .S(
        my_filter_data_sum[71]) );
  FA_X1 my_filter_adder_mult_4_addition_add_19_U1_2 ( .A(
        my_filter_adder_mult_4_res_mult[2]), .B(my_filter_data_sum[86]), .CI(
        my_filter_adder_mult_4_addition_add_19_carry[2]), .CO(
        my_filter_adder_mult_4_addition_add_19_carry[3]), .S(
        my_filter_data_sum[72]) );
  FA_X1 my_filter_adder_mult_4_addition_add_19_U1_3 ( .A(
        my_filter_adder_mult_4_res_mult[3]), .B(my_filter_data_sum[87]), .CI(
        my_filter_adder_mult_4_addition_add_19_carry[3]), .CO(
        my_filter_adder_mult_4_addition_add_19_carry[4]), .S(
        my_filter_data_sum[73]) );
  FA_X1 my_filter_adder_mult_4_addition_add_19_U1_4 ( .A(
        my_filter_adder_mult_4_res_mult[4]), .B(my_filter_data_sum[88]), .CI(
        my_filter_adder_mult_4_addition_add_19_carry[4]), .CO(
        my_filter_adder_mult_4_addition_add_19_carry[5]), .S(
        my_filter_data_sum[74]) );
  FA_X1 my_filter_adder_mult_4_addition_add_19_U1_5 ( .A(
        my_filter_adder_mult_4_res_mult[5]), .B(my_filter_data_sum[89]), .CI(
        my_filter_adder_mult_4_addition_add_19_carry[5]), .CO(
        my_filter_adder_mult_4_addition_add_19_carry[6]), .S(
        my_filter_data_sum[75]) );
  FA_X1 my_filter_adder_mult_4_addition_add_19_U1_6 ( .A(
        my_filter_adder_mult_4_res_mult[6]), .B(my_filter_data_sum[90]), .CI(
        my_filter_adder_mult_4_addition_add_19_carry[6]), .CO(
        my_filter_adder_mult_4_addition_add_19_carry[7]), .S(
        my_filter_data_sum[76]) );
  FA_X1 my_filter_adder_mult_4_addition_add_19_U1_7 ( .A(
        my_filter_adder_mult_4_res_mult[7]), .B(my_filter_data_sum[91]), .CI(
        my_filter_adder_mult_4_addition_add_19_carry[7]), .CO(
        my_filter_adder_mult_4_addition_add_19_carry[8]), .S(
        my_filter_data_sum[77]) );
  FA_X1 my_filter_adder_mult_4_addition_add_19_U1_8 ( .A(
        my_filter_adder_mult_4_res_mult[8]), .B(my_filter_data_sum[92]), .CI(
        my_filter_adder_mult_4_addition_add_19_carry[8]), .CO(
        my_filter_adder_mult_4_addition_add_19_carry[9]), .S(
        my_filter_data_sum[78]) );
  FA_X1 my_filter_adder_mult_4_addition_add_19_U1_9 ( .A(
        my_filter_adder_mult_4_res_mult[9]), .B(my_filter_data_sum[93]), .CI(
        my_filter_adder_mult_4_addition_add_19_carry[9]), .CO(
        my_filter_adder_mult_4_addition_add_19_carry[10]), .S(
        my_filter_data_sum[79]) );
  FA_X1 my_filter_adder_mult_4_addition_add_19_U1_10 ( .A(
        my_filter_adder_mult_4_res_mult[10]), .B(my_filter_data_sum[94]), .CI(
        my_filter_adder_mult_4_addition_add_19_carry[10]), .CO(
        my_filter_adder_mult_4_addition_add_19_carry[11]), .S(
        my_filter_data_sum[80]) );
  FA_X1 my_filter_adder_mult_4_addition_add_19_U1_11 ( .A(
        my_filter_adder_mult_4_res_mult[11]), .B(my_filter_data_sum[95]), .CI(
        my_filter_adder_mult_4_addition_add_19_carry[11]), .CO(
        my_filter_adder_mult_4_addition_add_19_carry[12]), .S(
        my_filter_data_sum[81]) );
  FA_X1 my_filter_adder_mult_4_addition_add_19_U1_12 ( .A(
        my_filter_adder_mult_4_res_mult[12]), .B(my_filter_data_sum[96]), .CI(
        my_filter_adder_mult_4_addition_add_19_carry[12]), .CO(
        my_filter_adder_mult_4_addition_add_19_carry[13]), .S(
        my_filter_data_sum[82]) );
  FA_X1 my_filter_adder_mult_4_addition_add_19_U1_13 ( .A(
        my_filter_adder_mult_4_res_mult[13]), .B(my_filter_data_sum[97]), .CI(
        my_filter_adder_mult_4_addition_add_19_carry[13]), .S(
        my_filter_data_sum[83]) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U276 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_12__12_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U275 ( .A1(
        my_filter_q_reg_chain_6__11_), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_11__13_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U274 ( .A1(
        my_filter_q_reg_coeff[67]), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_13__11_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U273 ( .A1(
        my_filter_q_reg_coeff[68]), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_13__12_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U272 ( .A1(
        my_filter_q_reg_chain_6__12_), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_12__13_) );
  INV_X1 my_filter_adder_mult_5_multiplication_mult_21_U271 ( .A(
        my_filter_q_reg_chain_6__12_), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_n87) );
  INV_X1 my_filter_adder_mult_5_multiplication_mult_21_U270 ( .A(
        my_filter_q_reg_chain_6__11_), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_n88) );
  INV_X1 my_filter_adder_mult_5_multiplication_mult_21_U269 ( .A(
        my_filter_q_reg_chain_6__13_), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_n86) );
  AND3_X1 my_filter_adder_mult_5_multiplication_mult_21_U268 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_ab_1__1_), .A2(
        my_filter_q_reg_coeff[56]), .A3(my_filter_q_reg_chain_6__0_), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_1__0_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U267 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_11__12_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U266 ( .A1(
        my_filter_q_reg_chain_6__10_), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_10__13_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U265 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_10__12_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U264 ( .A1(
        my_filter_q_reg_chain_6__9_), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_9__13_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U263 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n101), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_9__12_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U262 ( .A1(
        my_filter_q_reg_chain_6__8_), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_8__13_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U261 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_8__12_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U260 ( .A1(
        my_filter_q_reg_chain_6__7_), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_7__13_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U259 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_7__12_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U258 ( .A1(
        my_filter_q_reg_chain_6__6_), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_6__13_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U257 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_6__12_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U256 ( .A1(
        my_filter_q_reg_chain_6__5_), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_5__13_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U255 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_5__12_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U254 ( .A1(
        my_filter_q_reg_chain_6__4_), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_4__13_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U253 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_4__12_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U252 ( .A1(
        my_filter_q_reg_chain_6__3_), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_3__13_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U251 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_3__12_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U250 ( .A1(
        my_filter_q_reg_chain_6__2_), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_2__13_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U249 ( .A1(
        my_filter_q_reg_coeff[66]), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_13__10_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U248 ( .A1(
        my_filter_q_reg_coeff[64]), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_13__8_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U247 ( .A1(
        my_filter_q_reg_coeff[65]), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_13__9_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U246 ( .A1(
        my_filter_q_reg_coeff[62]), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_13__6_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U245 ( .A1(
        my_filter_q_reg_coeff[63]), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_13__7_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U244 ( .A1(
        my_filter_q_reg_coeff[60]), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_13__4_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U243 ( .A1(
        my_filter_q_reg_coeff[61]), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_13__5_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U242 ( .A1(
        my_filter_q_reg_coeff[59]), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_13__3_) );
  INV_X1 my_filter_adder_mult_5_multiplication_mult_21_U241 ( .A(
        my_filter_q_reg_coeff[56]), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_n113) );
  INV_X1 my_filter_adder_mult_5_multiplication_mult_21_U240 ( .A(
        my_filter_q_reg_coeff[57]), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_n112) );
  INV_X1 my_filter_adder_mult_5_multiplication_mult_21_U239 ( .A(
        my_filter_q_reg_chain_6__9_), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_n90) );
  INV_X1 my_filter_adder_mult_5_multiplication_mult_21_U238 ( .A(
        my_filter_q_reg_coeff[66]), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_n103) );
  INV_X1 my_filter_adder_mult_5_multiplication_mult_21_U237 ( .A(
        my_filter_q_reg_coeff[64]), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_n105) );
  INV_X1 my_filter_adder_mult_5_multiplication_mult_21_U236 ( .A(
        my_filter_q_reg_coeff[65]), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_n104) );
  INV_X1 my_filter_adder_mult_5_multiplication_mult_21_U235 ( .A(
        my_filter_q_reg_coeff[61]), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_n108) );
  INV_X1 my_filter_adder_mult_5_multiplication_mult_21_U234 ( .A(
        my_filter_q_reg_coeff[62]), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_n107) );
  INV_X1 my_filter_adder_mult_5_multiplication_mult_21_U233 ( .A(
        my_filter_q_reg_coeff[63]), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_n106) );
  INV_X1 my_filter_adder_mult_5_multiplication_mult_21_U232 ( .A(
        my_filter_q_reg_coeff[58]), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_n111) );
  INV_X1 my_filter_adder_mult_5_multiplication_mult_21_U231 ( .A(
        my_filter_q_reg_coeff[59]), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_n110) );
  INV_X1 my_filter_adder_mult_5_multiplication_mult_21_U230 ( .A(
        my_filter_q_reg_coeff[60]), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_n109) );
  INV_X1 my_filter_adder_mult_5_multiplication_mult_21_U229 ( .A(
        my_filter_q_reg_chain_6__10_), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_n89) );
  INV_X1 my_filter_adder_mult_5_multiplication_mult_21_U228 ( .A(
        my_filter_q_reg_chain_6__8_), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_n91) );
  INV_X1 my_filter_adder_mult_5_multiplication_mult_21_U227 ( .A(
        my_filter_q_reg_chain_6__7_), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_n92) );
  INV_X1 my_filter_adder_mult_5_multiplication_mult_21_U226 ( .A(
        my_filter_q_reg_chain_6__6_), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_n93) );
  INV_X1 my_filter_adder_mult_5_multiplication_mult_21_U225 ( .A(
        my_filter_q_reg_chain_6__5_), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_n94) );
  INV_X1 my_filter_adder_mult_5_multiplication_mult_21_U224 ( .A(
        my_filter_q_reg_chain_6__4_), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_n95) );
  INV_X1 my_filter_adder_mult_5_multiplication_mult_21_U223 ( .A(
        my_filter_q_reg_chain_6__2_), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_n97) );
  INV_X1 my_filter_adder_mult_5_multiplication_mult_21_U222 ( .A(
        my_filter_q_reg_chain_6__3_), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_n96) );
  AND2_X1 my_filter_adder_mult_5_multiplication_mult_21_U221 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_ab_0__13_), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_ab_1__12_), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_n15) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U220 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_2__12_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U219 ( .A1(
        my_filter_q_reg_chain_6__1_), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_1__13_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U218 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_12__0_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U217 ( .A1(
        my_filter_q_reg_coeff[56]), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_13__0_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U216 ( .A1(
        my_filter_q_reg_coeff[57]), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_13__1_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U215 ( .A1(
        my_filter_q_reg_coeff[58]), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_13__2_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U214 ( .A1(
        my_filter_q_reg_chain_6__0_), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_0__13_) );
  INV_X1 my_filter_adder_mult_5_multiplication_mult_21_U213 ( .A(
        my_filter_q_reg_coeff[69]), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_n100) );
  INV_X1 my_filter_adder_mult_5_multiplication_mult_21_U212 ( .A(
        my_filter_q_reg_chain_6__0_), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_n99) );
  INV_X1 my_filter_adder_mult_5_multiplication_mult_21_U211 ( .A(
        my_filter_q_reg_chain_6__1_), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_n98) );
  INV_X1 my_filter_adder_mult_5_multiplication_mult_21_U210 ( .A(
        my_filter_q_reg_coeff[68]), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_n101) );
  INV_X1 my_filter_adder_mult_5_multiplication_mult_21_U209 ( .A(
        my_filter_q_reg_coeff[67]), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_n102) );
  AND2_X1 my_filter_adder_mult_5_multiplication_mult_21_U208 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_13__12_), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_13__13_), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_n3) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U207 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n100), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_13__13_) );
  AND2_X1 my_filter_adder_mult_5_multiplication_mult_21_U206 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_13__9_), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_13__10_), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_n49) );
  AND2_X1 my_filter_adder_mult_5_multiplication_mult_21_U205 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_13__10_), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_13__11_), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_n51) );
  AND2_X1 my_filter_adder_mult_5_multiplication_mult_21_U204 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_13__7_), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_13__8_), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_n48) );
  AND2_X1 my_filter_adder_mult_5_multiplication_mult_21_U203 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_13__5_), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_13__6_), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_n47) );
  AND2_X1 my_filter_adder_mult_5_multiplication_mult_21_U202 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_13__3_), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_13__4_), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_n38) );
  AND2_X1 my_filter_adder_mult_5_multiplication_mult_21_U201 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_13__1_), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_13__2_), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_n46) );
  AND2_X1 my_filter_adder_mult_5_multiplication_mult_21_U200 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_13__8_), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_13__9_), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_n39) );
  AND2_X1 my_filter_adder_mult_5_multiplication_mult_21_U199 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_13__6_), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_13__7_), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_n44) );
  AND2_X1 my_filter_adder_mult_5_multiplication_mult_21_U198 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_13__4_), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_13__5_), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_n43) );
  AND2_X1 my_filter_adder_mult_5_multiplication_mult_21_U197 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_13__2_), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_13__3_), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_n42) );
  AND2_X1 my_filter_adder_mult_5_multiplication_mult_21_U196 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_13__0_), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_13__1_), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_n31) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U195 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_8__0_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U194 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n113), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_9__0_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U193 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_8__1_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U192 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_6__0_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U191 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_7__0_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U190 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_7__1_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U189 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_6__1_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U188 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_6__3_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U187 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_4__0_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U186 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_5__0_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U185 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_5__1_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U184 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_5__3_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U183 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_5__4_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U182 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_4__1_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U181 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_4__3_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U180 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_4__5_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U179 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_2__0_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U178 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_3__0_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U177 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_3__1_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U176 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_3__3_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U175 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_3__4_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U174 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_3__5_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U173 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_3__6_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U172 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_12__11_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U171 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_12__9_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U170 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_12__10_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U169 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_11__10_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U168 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_11__11_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U167 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_12__7_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U166 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_12__8_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U165 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_10__11_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U164 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_11__8_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U163 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_11__9_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U162 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_12__5_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U161 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_12__6_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U160 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_10__9_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U159 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_10__10_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U158 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_11__6_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U157 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_11__7_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U156 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n103), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_9__10_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U155 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n102), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_9__11_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U154 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_12__4_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U153 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_10__7_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U152 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_10__8_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U151 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_8__11_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U150 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_11__5_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U149 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n105), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_9__8_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U148 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n104), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_9__9_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U147 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_10__6_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U146 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_8__9_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U145 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_8__10_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U144 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n106), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_9__7_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U143 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_7__10_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U142 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_7__11_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U141 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_8__8_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U140 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_6__11_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U139 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_7__9_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U138 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_6__10_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U137 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_7__2_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U136 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_5__11_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U135 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_6__2_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U134 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_4__11_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U133 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_5__2_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U132 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_4__2_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U131 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_4__4_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U130 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_3__2_) );
  AND2_X1 my_filter_adder_mult_5_multiplication_mult_21_U129 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_ab_0__2_), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_ab_1__1_), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_n14) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U128 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_2__1_) );
  AND2_X1 my_filter_adder_mult_5_multiplication_mult_21_U127 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_ab_0__3_), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_ab_1__2_), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_n13) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U126 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_2__2_) );
  AND2_X1 my_filter_adder_mult_5_multiplication_mult_21_U125 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_ab_0__4_), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_ab_1__3_), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_n12) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U124 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_2__3_) );
  AND2_X1 my_filter_adder_mult_5_multiplication_mult_21_U123 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_ab_0__5_), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_ab_1__4_), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_n11) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U122 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_2__4_) );
  AND2_X1 my_filter_adder_mult_5_multiplication_mult_21_U121 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_ab_0__6_), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_ab_1__5_), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_n10) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U120 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_2__5_) );
  AND2_X1 my_filter_adder_mult_5_multiplication_mult_21_U119 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_ab_0__7_), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_ab_1__6_), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_n9) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U118 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_2__6_) );
  AND2_X1 my_filter_adder_mult_5_multiplication_mult_21_U117 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_ab_0__8_), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_ab_1__7_), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_n8) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U116 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_2__7_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U115 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_1__2_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U114 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_1__3_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U113 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_1__4_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U112 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_1__5_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U111 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_1__6_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U110 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_1__7_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U109 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_1__8_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U108 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_1__9_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U107 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_0__2_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U106 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_0__3_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U105 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_0__4_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U104 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_0__5_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U103 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_0__6_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U102 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_0__7_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U101 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_0__8_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U100 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_0__9_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U99 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n98), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n112), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_1__1_) );
  AND2_X1 my_filter_adder_mult_5_multiplication_mult_21_U98 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_13__11_), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_13__12_), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_n52) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U97 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_12__1_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U96 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_10__0_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U95 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_11__0_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U94 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_11__1_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U93 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_10__1_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U92 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n112), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_9__1_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U91 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n110), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_9__3_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U90 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_8__3_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U89 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_7__3_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U88 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_7__4_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U87 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_7__5_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U86 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_6__5_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U85 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_5__5_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U84 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_5__6_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U83 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_5__7_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U82 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_3__7_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U81 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_3__8_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U80 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_3__9_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U79 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_12__2_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U78 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_12__3_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U77 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_11__3_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U76 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_11__4_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U75 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_10__4_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U74 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_10__5_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U73 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_11__2_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U72 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n108), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_9__5_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U71 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n107), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_9__6_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U70 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_10__2_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U69 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_10__3_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U68 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_8__6_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U67 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_8__7_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U66 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n111), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_9__2_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U65 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n109), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_9__4_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U64 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_7__7_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U63 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_7__8_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U62 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_8__2_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U61 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_8__4_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U60 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_8__5_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U59 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_6__8_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U58 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_6__9_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U57 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_7__6_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U56 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_5__9_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U55 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_5__10_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U54 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_6__4_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U52 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_6__6_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U51 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_6__7_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U49 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_4__10_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U48 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_5__8_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U47 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_3__11_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U46 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_4__6_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U44 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_4__7_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U43 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_4__8_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U42 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_4__9_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U39 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_3__10_) );
  AND2_X1 my_filter_adder_mult_5_multiplication_mult_21_U38 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_ab_0__9_), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_ab_1__8_), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_n7) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U31 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_2__8_) );
  AND2_X1 my_filter_adder_mult_5_multiplication_mult_21_U14 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_ab_0__10_), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_ab_1__9_), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_n6) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U13 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_2__9_) );
  AND2_X1 my_filter_adder_mult_5_multiplication_mult_21_U12 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_ab_0__11_), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_ab_1__10_), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_n5) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U11 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_2__10_) );
  AND2_X1 my_filter_adder_mult_5_multiplication_mult_21_U10 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_ab_0__12_), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_ab_1__11_), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_n4) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U9 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_2__11_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U8 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_1__12_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U7 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_1__10_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U6 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_1__11_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U5 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_0__10_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U4 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_0__11_) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U3 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_ab_0__12_) );
  INV_X1 my_filter_adder_mult_5_multiplication_mult_21_U2 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_13__13_), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_n85) );
  XOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U50 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_13__11_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_13__12_), .Z(
        my_filter_adder_mult_5_multiplication_mult_21_n50) );
  XOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U45 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_13__10_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_13__11_), .Z(
        my_filter_adder_mult_5_multiplication_mult_21_n45) );
  XOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U41 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_13__5_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_13__6_), .Z(
        my_filter_adder_mult_5_multiplication_mult_21_n41) );
  XOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U40 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_13__3_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_13__4_), .Z(
        my_filter_adder_mult_5_multiplication_mult_21_n40) );
  XOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U37 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_13__8_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_13__9_), .Z(
        my_filter_adder_mult_5_multiplication_mult_21_n37) );
  XOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U36 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_13__9_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_13__10_), .Z(
        my_filter_adder_mult_5_multiplication_mult_21_n36) );
  XOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U35 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_13__6_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_13__7_), .Z(
        my_filter_adder_mult_5_multiplication_mult_21_n35) );
  XOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U34 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_13__7_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_13__8_), .Z(
        my_filter_adder_mult_5_multiplication_mult_21_n34) );
  XOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U33 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_13__4_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_13__5_), .Z(
        my_filter_adder_mult_5_multiplication_mult_21_n33) );
  XOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U32 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_13__2_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_13__3_), .Z(
        my_filter_adder_mult_5_multiplication_mult_21_n32) );
  XOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U30 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_13__1_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_13__2_), .Z(
        my_filter_adder_mult_5_multiplication_mult_21_n30) );
  XOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U29 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_13__0_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_13__1_), .Z(
        my_filter_adder_mult_5_multiplication_mult_21_n29) );
  XOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U27 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_1__1_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_ab_0__2_), .Z(
        my_filter_adder_mult_5_multiplication_mult_21_n28) );
  XOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U26 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_13__12_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_13__13_), .Z(
        my_filter_adder_mult_5_multiplication_mult_21_n27) );
  XOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U25 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_1__12_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_ab_0__13_), .Z(
        my_filter_adder_mult_5_multiplication_mult_21_n26) );
  XOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U24 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_1__2_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_ab_0__3_), .Z(
        my_filter_adder_mult_5_multiplication_mult_21_n25) );
  XOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U23 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_1__3_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_ab_0__4_), .Z(
        my_filter_adder_mult_5_multiplication_mult_21_n24) );
  XOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U22 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_1__4_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_ab_0__5_), .Z(
        my_filter_adder_mult_5_multiplication_mult_21_n23) );
  XOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U21 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_1__5_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_ab_0__6_), .Z(
        my_filter_adder_mult_5_multiplication_mult_21_n22) );
  XOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U20 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_1__6_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_ab_0__7_), .Z(
        my_filter_adder_mult_5_multiplication_mult_21_n21) );
  XOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U19 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_1__7_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_ab_0__8_), .Z(
        my_filter_adder_mult_5_multiplication_mult_21_n20) );
  XOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U18 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_1__8_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_ab_0__9_), .Z(
        my_filter_adder_mult_5_multiplication_mult_21_n19) );
  XOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U17 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_1__9_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_ab_0__10_), .Z(
        my_filter_adder_mult_5_multiplication_mult_21_n18) );
  XOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U16 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_1__10_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_ab_0__11_), .Z(
        my_filter_adder_mult_5_multiplication_mult_21_n17) );
  XOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_U15 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_1__11_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_ab_0__12_), .Z(
        my_filter_adder_mult_5_multiplication_mult_21_n16) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S3_2_12 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_2__12_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_n15), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_ab_1__13_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_2__12_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_2__12_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_2_11 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_2__11_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_n4), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_n26), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_2__11_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_2__11_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_2_10 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_2__10_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_n5), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_n16), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_2__10_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_2__10_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_2_9 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_2__9_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_n6), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_n17), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_2__9_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_2__9_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_2_8 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_2__8_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_n7), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_n18), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_2__8_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_2__8_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_2_7 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_2__7_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_n8), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_n19), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_2__7_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_2__7_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_2_6 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_2__6_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_n9), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_n20), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_2__6_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_2__6_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_2_5 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_2__5_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_n10), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_n21), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_2__5_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_2__5_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_2_4 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_2__4_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_n11), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_n22), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_2__4_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_2__4_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_2_3 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_2__3_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_n12), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_n23), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_2__3_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_2__3_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_2_2 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_2__2_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_n13), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_n24), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_2__2_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_2__2_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_2_1 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_2__1_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_n14), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_n25), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_2__1_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_2__1_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S1_2_0 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_2__0_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_1__0_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_n28), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_2__0_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_A1_0_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S3_3_12 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_3__12_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_2__12_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_ab_2__13_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_3__12_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_3__12_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_3_11 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_3__11_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_2__11_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_2__12_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_3__11_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_3__11_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_3_10 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_3__10_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_2__10_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_2__11_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_3__10_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_3__10_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_3_9 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_3__9_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_2__9_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_2__10_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_3__9_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_3__9_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_3_8 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_3__8_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_2__8_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_2__9_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_3__8_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_3__8_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_3_7 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_3__7_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_2__7_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_2__8_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_3__7_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_3__7_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_3_6 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_3__6_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_2__6_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_2__7_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_3__6_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_3__6_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_3_5 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_3__5_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_2__5_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_2__6_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_3__5_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_3__5_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_3_4 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_3__4_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_2__4_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_2__5_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_3__4_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_3__4_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_3_3 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_3__3_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_2__3_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_2__4_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_3__3_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_3__3_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_3_2 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_3__2_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_2__2_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_2__3_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_3__2_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_3__2_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_3_1 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_3__1_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_2__1_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_2__2_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_3__1_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_3__1_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S1_3_0 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_3__0_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_2__0_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_2__1_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_3__0_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_A1_1_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S3_4_12 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_4__12_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_3__12_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_ab_3__13_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_4__12_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_4__12_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_4_11 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_4__11_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_3__11_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_3__12_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_4__11_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_4__11_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_4_10 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_4__10_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_3__10_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_3__11_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_4__10_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_4__10_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_4_9 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_4__9_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_3__9_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_3__10_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_4__9_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_4__9_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_4_8 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_4__8_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_3__8_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_3__9_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_4__8_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_4__8_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_4_7 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_4__7_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_3__7_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_3__8_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_4__7_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_4__7_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_4_6 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_4__6_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_3__6_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_3__7_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_4__6_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_4__6_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_4_5 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_4__5_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_3__5_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_3__6_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_4__5_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_4__5_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_4_4 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_4__4_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_3__4_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_3__5_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_4__4_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_4__4_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_4_3 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_4__3_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_3__3_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_3__4_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_4__3_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_4__3_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_4_2 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_4__2_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_3__2_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_3__3_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_4__2_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_4__2_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_4_1 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_4__1_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_3__1_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_3__2_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_4__1_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_4__1_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S1_4_0 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_4__0_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_3__0_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_3__1_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_4__0_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_A1_2_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S3_5_12 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_5__12_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_4__12_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_ab_4__13_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_5__12_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_5__12_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_5_11 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_5__11_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_4__11_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_4__12_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_5__11_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_5__11_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_5_10 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_5__10_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_4__10_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_4__11_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_5__10_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_5__10_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_5_9 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_5__9_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_4__9_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_4__10_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_5__9_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_5__9_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_5_8 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_5__8_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_4__8_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_4__9_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_5__8_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_5__8_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_5_7 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_5__7_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_4__7_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_4__8_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_5__7_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_5__7_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_5_6 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_5__6_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_4__6_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_4__7_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_5__6_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_5__6_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_5_5 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_5__5_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_4__5_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_4__6_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_5__5_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_5__5_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_5_4 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_5__4_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_4__4_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_4__5_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_5__4_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_5__4_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_5_3 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_5__3_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_4__3_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_4__4_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_5__3_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_5__3_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_5_2 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_5__2_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_4__2_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_4__3_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_5__2_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_5__2_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_5_1 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_5__1_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_4__1_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_4__2_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_5__1_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_5__1_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S1_5_0 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_5__0_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_4__0_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_4__1_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_5__0_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_A1_3_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S3_6_12 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_6__12_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_5__12_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_ab_5__13_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_6__12_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_6__12_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_6_11 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_6__11_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_5__11_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_5__12_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_6__11_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_6__11_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_6_10 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_6__10_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_5__10_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_5__11_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_6__10_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_6__10_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_6_9 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_6__9_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_5__9_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_5__10_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_6__9_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_6__9_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_6_8 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_6__8_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_5__8_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_5__9_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_6__8_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_6__8_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_6_7 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_6__7_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_5__7_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_5__8_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_6__7_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_6__7_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_6_6 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_6__6_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_5__6_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_5__7_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_6__6_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_6__6_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_6_5 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_6__5_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_5__5_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_5__6_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_6__5_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_6__5_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_6_4 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_6__4_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_5__4_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_5__5_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_6__4_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_6__4_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_6_3 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_6__3_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_5__3_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_5__4_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_6__3_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_6__3_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_6_2 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_6__2_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_5__2_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_5__3_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_6__2_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_6__2_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_6_1 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_6__1_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_5__1_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_5__2_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_6__1_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_6__1_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S1_6_0 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_6__0_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_5__0_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_5__1_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_6__0_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_A1_4_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S3_7_12 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_7__12_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_6__12_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_ab_6__13_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_7__12_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_7__12_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_7_11 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_7__11_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_6__11_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_6__12_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_7__11_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_7__11_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_7_10 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_7__10_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_6__10_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_6__11_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_7__10_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_7__10_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_7_9 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_7__9_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_6__9_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_6__10_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_7__9_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_7__9_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_7_8 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_7__8_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_6__8_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_6__9_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_7__8_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_7__8_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_7_7 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_7__7_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_6__7_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_6__8_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_7__7_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_7__7_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_7_6 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_7__6_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_6__6_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_6__7_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_7__6_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_7__6_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_7_5 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_7__5_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_6__5_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_6__6_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_7__5_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_7__5_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_7_4 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_7__4_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_6__4_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_6__5_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_7__4_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_7__4_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_7_3 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_7__3_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_6__3_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_6__4_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_7__3_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_7__3_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_7_2 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_7__2_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_6__2_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_6__3_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_7__2_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_7__2_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_7_1 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_7__1_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_6__1_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_6__2_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_7__1_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_7__1_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S1_7_0 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_7__0_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_6__0_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_6__1_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_7__0_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_A1_5_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S3_8_12 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_8__12_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_7__12_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_ab_7__13_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_8__12_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_8__12_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_8_11 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_8__11_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_7__11_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_7__12_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_8__11_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_8__11_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_8_10 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_8__10_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_7__10_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_7__11_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_8__10_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_8__10_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_8_9 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_8__9_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_7__9_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_7__10_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_8__9_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_8__9_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_8_8 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_8__8_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_7__8_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_7__9_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_8__8_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_8__8_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_8_7 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_8__7_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_7__7_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_7__8_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_8__7_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_8__7_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_8_6 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_8__6_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_7__6_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_7__7_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_8__6_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_8__6_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_8_5 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_8__5_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_7__5_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_7__6_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_8__5_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_8__5_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_8_4 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_8__4_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_7__4_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_7__5_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_8__4_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_8__4_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_8_3 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_8__3_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_7__3_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_7__4_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_8__3_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_8__3_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_8_2 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_8__2_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_7__2_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_7__3_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_8__2_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_8__2_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_8_1 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_8__1_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_7__1_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_7__2_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_8__1_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_8__1_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S1_8_0 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_8__0_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_7__0_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_7__1_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_8__0_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_A1_6_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S3_9_12 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_9__12_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_8__12_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_ab_8__13_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_9__12_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_9__12_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_9_11 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_9__11_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_8__11_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_8__12_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_9__11_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_9__11_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_9_10 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_9__10_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_8__10_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_8__11_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_9__10_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_9__10_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_9_9 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_9__9_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_8__9_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_8__10_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_9__9_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_9__9_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_9_8 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_9__8_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_8__8_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_8__9_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_9__8_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_9__8_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_9_7 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_9__7_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_8__7_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_8__8_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_9__7_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_9__7_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_9_6 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_9__6_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_8__6_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_8__7_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_9__6_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_9__6_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_9_5 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_9__5_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_8__5_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_8__6_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_9__5_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_9__5_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_9_4 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_9__4_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_8__4_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_8__5_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_9__4_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_9__4_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_9_3 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_9__3_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_8__3_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_8__4_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_9__3_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_9__3_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_9_2 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_9__2_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_8__2_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_8__3_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_9__2_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_9__2_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_9_1 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_9__1_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_8__1_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_8__2_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_9__1_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_9__1_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S1_9_0 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_9__0_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_8__0_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_8__1_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_9__0_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_A1_7_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S3_10_12 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_10__12_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_9__12_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_ab_9__13_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_10__12_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_10__12_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_10_11 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_10__11_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_9__11_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_9__12_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_10__11_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_10__11_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_10_10 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_10__10_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_9__10_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_9__11_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_10__10_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_10__10_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_10_9 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_10__9_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_9__9_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_9__10_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_10__9_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_10__9_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_10_8 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_10__8_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_9__8_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_9__9_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_10__8_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_10__8_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_10_7 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_10__7_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_9__7_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_9__8_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_10__7_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_10__7_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_10_6 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_10__6_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_9__6_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_9__7_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_10__6_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_10__6_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_10_5 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_10__5_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_9__5_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_9__6_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_10__5_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_10__5_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_10_4 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_10__4_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_9__4_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_9__5_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_10__4_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_10__4_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_10_3 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_10__3_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_9__3_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_9__4_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_10__3_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_10__3_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_10_2 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_10__2_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_9__2_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_9__3_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_10__2_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_10__2_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_10_1 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_10__1_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_9__1_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_9__2_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_10__1_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_10__1_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S1_10_0 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_10__0_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_9__0_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_9__1_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_10__0_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_A1_8_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S3_11_12 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_11__12_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_10__12_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_ab_10__13_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_11__12_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_11__12_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_11_11 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_11__11_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_10__11_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_10__12_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_11__11_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_11__11_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_11_10 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_11__10_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_10__10_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_10__11_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_11__10_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_11__10_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_11_9 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_11__9_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_10__9_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_10__10_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_11__9_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_11__9_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_11_8 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_11__8_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_10__8_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_10__9_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_11__8_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_11__8_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_11_7 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_11__7_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_10__7_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_10__8_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_11__7_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_11__7_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_11_6 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_11__6_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_10__6_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_10__7_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_11__6_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_11__6_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_11_5 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_11__5_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_10__5_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_10__6_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_11__5_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_11__5_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_11_4 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_11__4_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_10__4_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_10__5_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_11__4_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_11__4_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_11_3 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_11__3_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_10__3_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_10__4_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_11__3_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_11__3_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_11_2 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_11__2_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_10__2_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_10__3_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_11__2_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_11__2_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_11_1 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_11__1_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_10__1_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_10__2_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_11__1_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_11__1_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S1_11_0 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_11__0_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_10__0_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_10__1_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_11__0_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_A1_9_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S3_12_12 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_12__12_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_11__12_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_ab_11__13_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_12__12_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_12__12_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_12_11 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_12__11_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_11__11_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_11__12_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_12__11_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_12__11_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_12_10 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_12__10_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_11__10_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_11__11_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_12__10_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_12__10_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_12_9 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_12__9_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_11__9_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_11__10_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_12__9_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_12__9_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_12_8 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_12__8_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_11__8_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_11__9_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_12__8_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_12__8_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_12_7 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_12__7_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_11__7_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_11__8_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_12__7_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_12__7_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_12_6 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_12__6_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_11__6_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_11__7_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_12__6_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_12__6_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_12_5 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_12__5_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_11__5_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_11__6_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_12__5_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_12__5_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_12_4 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_12__4_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_11__4_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_11__5_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_12__4_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_12__4_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_12_3 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_12__3_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_11__3_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_11__4_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_12__3_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_12__3_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_12_2 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_12__2_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_11__2_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_11__3_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_12__2_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_12__2_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S2_12_1 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_12__1_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_11__1_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_11__2_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_12__1_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_12__1_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S1_12_0 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_12__0_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_11__0_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_11__1_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_12__0_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_A1_10_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S14_13 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_n86), .B(
        my_filter_adder_mult_5_multiplication_mult_21_n100), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_ab_13__13_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_13__13_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_13__13_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S5_12 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_13__12_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_12__12_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_ab_12__13_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_13__12_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_13__12_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S4_11 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_13__11_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_12__11_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_12__12_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_13__11_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_13__11_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S4_10 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_13__10_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_12__10_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_12__11_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_13__10_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_13__10_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S4_9 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_13__9_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_12__9_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_12__10_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_13__9_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_13__9_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S4_8 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_13__8_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_12__8_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_12__9_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_13__8_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_13__8_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S4_7 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_13__7_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_12__7_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_12__8_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_13__7_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_13__7_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S4_6 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_13__6_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_12__6_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_12__7_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_13__6_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_13__6_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S4_5 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_13__5_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_12__5_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_12__6_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_13__5_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_13__5_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S4_4 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_13__4_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_12__4_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_12__5_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_13__4_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_13__4_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S4_3 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_13__3_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_12__3_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_12__4_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_13__3_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_13__3_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S4_2 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_13__2_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_12__2_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_12__3_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_13__2_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_13__2_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S4_1 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_13__1_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_12__1_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_12__2_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_13__1_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_13__1_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S4_0 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_ab_13__0_), .B(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_12__0_), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_12__1_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_CARRYB_13__0_), .S(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_13__0_) );
  FA_X1 my_filter_adder_mult_5_multiplication_mult_21_S14_13_0 ( .A(
        my_filter_q_reg_chain_6__13_), .B(my_filter_q_reg_coeff[69]), .CI(
        my_filter_adder_mult_5_multiplication_mult_21_SUMB_13__0_), .CO(
        my_filter_adder_mult_5_multiplication_mult_21_A2_12_), .S(
        my_filter_adder_mult_5_res_mult[0]) );
  OAI21_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U72 ( .B1(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n15), .B2(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n16), .A(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n17), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n13) );
  NAND2_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U71 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_A2_12_), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n29), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n56) );
  OAI21_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U70 ( .B1(
        my_filter_adder_mult_5_multiplication_mult_21_A2_12_), .B2(
        my_filter_adder_mult_5_multiplication_mult_21_n29), .A(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n56), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n59) );
  INV_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U69 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n59), .ZN(
        my_filter_adder_mult_5_res_mult[1]) );
  AND2_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U68 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n49), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n45), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n20) );
  NAND2_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U66 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n51), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n50), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n17) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U65 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n51), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n50), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n15) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U64 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n49), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n45), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n21) );
  AND2_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U63 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n48), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n37), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n28) );
  AND2_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U61 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n47), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n35), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n36) );
  AND2_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U60 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n38), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n33), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n44) );
  AND2_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U59 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n46), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n32), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n52) );
  NAND2_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U58 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n39), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n36), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n25) );
  NAND2_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U56 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n44), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n34), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n33) );
  NAND2_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U55 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n43), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n41), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n41) );
  NAND2_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U54 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n42), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n40), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n49) );
  NAND2_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U53 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n31), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n30), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n57) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U51 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n39), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n36), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n23) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U50 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n44), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n34), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n31) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U49 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n43), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n41), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n39) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U48 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n42), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n40), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n47) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U46 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n48), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n37), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n29) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U45 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n47), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n35), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n37) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U44 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n38), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n33), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n45) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U43 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n46), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n32), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n53) );
  OAI21_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U41 ( .B1(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n55), .B2(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n56), .A(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n57), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n51) );
  INV_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U40 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n55), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n60) );
  NAND2_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U39 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n60), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n57), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n58) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U38 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_n31), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_n30), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n55) );
  OAI21_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U36 ( .B1(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n23), .B2(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n24), .A(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n25), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n19) );
  OAI21_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U35 ( .B1(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n31), .B2(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n32), .A(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n33), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n27) );
  OAI21_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U34 ( .B1(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n39), .B2(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n40), .A(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n41), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n35) );
  OAI21_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U33 ( .B1(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n47), .B2(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n48), .A(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n49), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n43) );
  INV_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U31 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n21), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n63) );
  AOI21_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U30 ( .B1(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n63), .B2(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n19), .A(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n20), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n16) );
  INV_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U29 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n29), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n71) );
  AOI21_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U28 ( .B1(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n71), .B2(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n27), .A(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n28), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n24) );
  INV_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U26 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n37), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n69) );
  AOI21_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U25 ( .B1(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n69), .B2(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n35), .A(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n36), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n32) );
  INV_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U24 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n45), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n67) );
  AOI21_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U23 ( .B1(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n67), .B2(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n43), .A(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n44), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n40) );
  INV_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U21 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n53), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n65) );
  AOI21_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U20 ( .B1(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n65), .B2(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n51), .A(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n52), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n48) );
  INV_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U19 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n15), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n62) );
  NAND2_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U18 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n62), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n17), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n18) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U16 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n20), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n21), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n22) );
  INV_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U13 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n23), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n64) );
  NAND2_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U12 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n64), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n25), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n26) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U11 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n28), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n29), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n30) );
  INV_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U10 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n31), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n70) );
  NAND2_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U9 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n70), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n33), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n34) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U8 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n36), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n37), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n38) );
  INV_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U7 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n39), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n68) );
  NAND2_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U6 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n68), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n41), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n42) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U5 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n44), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n45), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n46) );
  INV_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U4 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n47), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n66) );
  NAND2_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U3 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n66), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n49), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n50) );
  NOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U2 ( .A1(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n52), .A2(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n53), .ZN(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n54) );
  XOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U67 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n56), .B(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n58), .Z(
        my_filter_adder_mult_5_res_mult[2]) );
  XOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U62 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n51), .B(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n54), .Z(
        my_filter_adder_mult_5_res_mult[3]) );
  XOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U57 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n50), .B(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n48), .Z(
        my_filter_adder_mult_5_res_mult[4]) );
  XOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U52 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n43), .B(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n46), .Z(
        my_filter_adder_mult_5_res_mult[5]) );
  XOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U47 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n42), .B(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n40), .Z(
        my_filter_adder_mult_5_res_mult[6]) );
  XOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U42 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n35), .B(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n38), .Z(
        my_filter_adder_mult_5_res_mult[7]) );
  XOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U37 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n34), .B(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n32), .Z(
        my_filter_adder_mult_5_res_mult[8]) );
  XOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U32 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n27), .B(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n30), .Z(
        my_filter_adder_mult_5_res_mult[9]) );
  XOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U27 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n26), .B(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n24), .Z(
        my_filter_adder_mult_5_res_mult[10]) );
  XOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U22 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n19), .B(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n22), .Z(
        my_filter_adder_mult_5_res_mult[11]) );
  XOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U17 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n18), .B(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n16), .Z(
        my_filter_adder_mult_5_res_mult[12]) );
  XOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U15 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_n52), .B(
        my_filter_adder_mult_5_multiplication_mult_21_n27), .Z(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n14) );
  XOR2_X1 my_filter_adder_mult_5_multiplication_mult_21_FS_1_U14 ( .A(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n13), .B(
        my_filter_adder_mult_5_multiplication_mult_21_FS_1_n14), .Z(
        my_filter_adder_mult_5_res_mult[13]) );
  AND2_X1 my_filter_adder_mult_5_addition_add_19_U1 ( .A1(
        my_filter_data_sum[70]), .A2(my_filter_adder_mult_5_res_mult[0]), .ZN(
        my_filter_adder_mult_5_addition_add_19_n1) );
  XOR2_X1 my_filter_adder_mult_5_addition_add_19_U2 ( .A(
        my_filter_data_sum[70]), .B(my_filter_adder_mult_5_res_mult[0]), .Z(
        my_filter_data_sum[56]) );
  FA_X1 my_filter_adder_mult_5_addition_add_19_U1_1 ( .A(
        my_filter_adder_mult_5_res_mult[1]), .B(my_filter_data_sum[71]), .CI(
        my_filter_adder_mult_5_addition_add_19_n1), .CO(
        my_filter_adder_mult_5_addition_add_19_carry[2]), .S(
        my_filter_data_sum[57]) );
  FA_X1 my_filter_adder_mult_5_addition_add_19_U1_2 ( .A(
        my_filter_adder_mult_5_res_mult[2]), .B(my_filter_data_sum[72]), .CI(
        my_filter_adder_mult_5_addition_add_19_carry[2]), .CO(
        my_filter_adder_mult_5_addition_add_19_carry[3]), .S(
        my_filter_data_sum[58]) );
  FA_X1 my_filter_adder_mult_5_addition_add_19_U1_3 ( .A(
        my_filter_adder_mult_5_res_mult[3]), .B(my_filter_data_sum[73]), .CI(
        my_filter_adder_mult_5_addition_add_19_carry[3]), .CO(
        my_filter_adder_mult_5_addition_add_19_carry[4]), .S(
        my_filter_data_sum[59]) );
  FA_X1 my_filter_adder_mult_5_addition_add_19_U1_4 ( .A(
        my_filter_adder_mult_5_res_mult[4]), .B(my_filter_data_sum[74]), .CI(
        my_filter_adder_mult_5_addition_add_19_carry[4]), .CO(
        my_filter_adder_mult_5_addition_add_19_carry[5]), .S(
        my_filter_data_sum[60]) );
  FA_X1 my_filter_adder_mult_5_addition_add_19_U1_5 ( .A(
        my_filter_adder_mult_5_res_mult[5]), .B(my_filter_data_sum[75]), .CI(
        my_filter_adder_mult_5_addition_add_19_carry[5]), .CO(
        my_filter_adder_mult_5_addition_add_19_carry[6]), .S(
        my_filter_data_sum[61]) );
  FA_X1 my_filter_adder_mult_5_addition_add_19_U1_6 ( .A(
        my_filter_adder_mult_5_res_mult[6]), .B(my_filter_data_sum[76]), .CI(
        my_filter_adder_mult_5_addition_add_19_carry[6]), .CO(
        my_filter_adder_mult_5_addition_add_19_carry[7]), .S(
        my_filter_data_sum[62]) );
  FA_X1 my_filter_adder_mult_5_addition_add_19_U1_7 ( .A(
        my_filter_adder_mult_5_res_mult[7]), .B(my_filter_data_sum[77]), .CI(
        my_filter_adder_mult_5_addition_add_19_carry[7]), .CO(
        my_filter_adder_mult_5_addition_add_19_carry[8]), .S(
        my_filter_data_sum[63]) );
  FA_X1 my_filter_adder_mult_5_addition_add_19_U1_8 ( .A(
        my_filter_adder_mult_5_res_mult[8]), .B(my_filter_data_sum[78]), .CI(
        my_filter_adder_mult_5_addition_add_19_carry[8]), .CO(
        my_filter_adder_mult_5_addition_add_19_carry[9]), .S(
        my_filter_data_sum[64]) );
  FA_X1 my_filter_adder_mult_5_addition_add_19_U1_9 ( .A(
        my_filter_adder_mult_5_res_mult[9]), .B(my_filter_data_sum[79]), .CI(
        my_filter_adder_mult_5_addition_add_19_carry[9]), .CO(
        my_filter_adder_mult_5_addition_add_19_carry[10]), .S(
        my_filter_data_sum[65]) );
  FA_X1 my_filter_adder_mult_5_addition_add_19_U1_10 ( .A(
        my_filter_adder_mult_5_res_mult[10]), .B(my_filter_data_sum[80]), .CI(
        my_filter_adder_mult_5_addition_add_19_carry[10]), .CO(
        my_filter_adder_mult_5_addition_add_19_carry[11]), .S(
        my_filter_data_sum[66]) );
  FA_X1 my_filter_adder_mult_5_addition_add_19_U1_11 ( .A(
        my_filter_adder_mult_5_res_mult[11]), .B(my_filter_data_sum[81]), .CI(
        my_filter_adder_mult_5_addition_add_19_carry[11]), .CO(
        my_filter_adder_mult_5_addition_add_19_carry[12]), .S(
        my_filter_data_sum[67]) );
  FA_X1 my_filter_adder_mult_5_addition_add_19_U1_12 ( .A(
        my_filter_adder_mult_5_res_mult[12]), .B(my_filter_data_sum[82]), .CI(
        my_filter_adder_mult_5_addition_add_19_carry[12]), .CO(
        my_filter_adder_mult_5_addition_add_19_carry[13]), .S(
        my_filter_data_sum[68]) );
  FA_X1 my_filter_adder_mult_5_addition_add_19_U1_13 ( .A(
        my_filter_adder_mult_5_res_mult[13]), .B(my_filter_data_sum[83]), .CI(
        my_filter_adder_mult_5_addition_add_19_carry[13]), .S(
        my_filter_data_sum[69]) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U276 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_12__12_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U275 ( .A1(
        my_filter_q_reg_chain_7__11_), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_11__13_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U274 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_11__12_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U273 ( .A1(
        my_filter_q_reg_chain_7__10_), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_10__13_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U272 ( .A1(
        my_filter_q_reg_coeff[52]), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_13__10_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U271 ( .A1(
        my_filter_q_reg_coeff[53]), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_13__11_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U270 ( .A1(
        my_filter_q_reg_coeff[54]), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_13__12_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U269 ( .A1(
        my_filter_q_reg_chain_7__12_), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_12__13_) );
  INV_X1 my_filter_adder_mult_6_multiplication_mult_21_U268 ( .A(
        my_filter_q_reg_chain_7__9_), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_n90) );
  INV_X1 my_filter_adder_mult_6_multiplication_mult_21_U267 ( .A(
        my_filter_q_reg_chain_7__12_), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_n87) );
  INV_X1 my_filter_adder_mult_6_multiplication_mult_21_U266 ( .A(
        my_filter_q_reg_chain_7__11_), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_n88) );
  INV_X1 my_filter_adder_mult_6_multiplication_mult_21_U265 ( .A(
        my_filter_q_reg_chain_7__10_), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_n89) );
  INV_X1 my_filter_adder_mult_6_multiplication_mult_21_U264 ( .A(
        my_filter_q_reg_chain_7__13_), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_n86) );
  AND2_X1 my_filter_adder_mult_6_multiplication_mult_21_U263 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_ab_0__13_), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_ab_1__12_), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_n15) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U262 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_2__12_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U261 ( .A1(
        my_filter_q_reg_chain_7__1_), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_1__13_) );
  AND3_X1 my_filter_adder_mult_6_multiplication_mult_21_U260 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_ab_1__1_), .A2(
        my_filter_q_reg_coeff[42]), .A3(my_filter_q_reg_chain_7__0_), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_1__0_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U259 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_12__0_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U258 ( .A1(
        my_filter_q_reg_coeff[42]), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_13__0_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U257 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_10__12_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U256 ( .A1(
        my_filter_q_reg_chain_7__9_), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_9__13_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U255 ( .A1(
        my_filter_q_reg_chain_7__8_), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_8__13_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U254 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n101), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_9__12_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U253 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_8__12_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U252 ( .A1(
        my_filter_q_reg_chain_7__7_), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_7__13_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U251 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_7__12_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U250 ( .A1(
        my_filter_q_reg_chain_7__6_), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_6__13_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U249 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_6__12_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U248 ( .A1(
        my_filter_q_reg_chain_7__5_), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_5__13_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U247 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_5__12_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U246 ( .A1(
        my_filter_q_reg_chain_7__4_), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_4__13_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U245 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_4__12_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U244 ( .A1(
        my_filter_q_reg_chain_7__3_), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_3__13_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U243 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_3__12_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U242 ( .A1(
        my_filter_q_reg_chain_7__2_), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_2__13_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U241 ( .A1(
        my_filter_q_reg_coeff[50]), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_13__8_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U240 ( .A1(
        my_filter_q_reg_coeff[51]), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_13__9_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U239 ( .A1(
        my_filter_q_reg_coeff[48]), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_13__6_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U238 ( .A1(
        my_filter_q_reg_coeff[49]), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_13__7_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U237 ( .A1(
        my_filter_q_reg_coeff[46]), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_13__4_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U236 ( .A1(
        my_filter_q_reg_coeff[47]), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_13__5_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U235 ( .A1(
        my_filter_q_reg_coeff[43]), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_13__1_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U234 ( .A1(
        my_filter_q_reg_coeff[44]), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_13__2_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U233 ( .A1(
        my_filter_q_reg_coeff[45]), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_13__3_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U232 ( .A1(
        my_filter_q_reg_chain_7__0_), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_0__13_) );
  INV_X1 my_filter_adder_mult_6_multiplication_mult_21_U231 ( .A(
        my_filter_q_reg_coeff[55]), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_n100) );
  INV_X1 my_filter_adder_mult_6_multiplication_mult_21_U230 ( .A(
        my_filter_q_reg_coeff[42]), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_n113) );
  INV_X1 my_filter_adder_mult_6_multiplication_mult_21_U229 ( .A(
        my_filter_q_reg_chain_7__0_), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_n99) );
  INV_X1 my_filter_adder_mult_6_multiplication_mult_21_U228 ( .A(
        my_filter_q_reg_coeff[43]), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_n112) );
  INV_X1 my_filter_adder_mult_6_multiplication_mult_21_U227 ( .A(
        my_filter_q_reg_chain_7__1_), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_n98) );
  INV_X1 my_filter_adder_mult_6_multiplication_mult_21_U226 ( .A(
        my_filter_q_reg_coeff[54]), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_n101) );
  INV_X1 my_filter_adder_mult_6_multiplication_mult_21_U225 ( .A(
        my_filter_q_reg_coeff[52]), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_n103) );
  INV_X1 my_filter_adder_mult_6_multiplication_mult_21_U224 ( .A(
        my_filter_q_reg_coeff[53]), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_n102) );
  INV_X1 my_filter_adder_mult_6_multiplication_mult_21_U223 ( .A(
        my_filter_q_reg_coeff[50]), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_n105) );
  INV_X1 my_filter_adder_mult_6_multiplication_mult_21_U222 ( .A(
        my_filter_q_reg_coeff[51]), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_n104) );
  INV_X1 my_filter_adder_mult_6_multiplication_mult_21_U221 ( .A(
        my_filter_q_reg_coeff[47]), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_n108) );
  INV_X1 my_filter_adder_mult_6_multiplication_mult_21_U220 ( .A(
        my_filter_q_reg_coeff[48]), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_n107) );
  INV_X1 my_filter_adder_mult_6_multiplication_mult_21_U219 ( .A(
        my_filter_q_reg_coeff[49]), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_n106) );
  INV_X1 my_filter_adder_mult_6_multiplication_mult_21_U218 ( .A(
        my_filter_q_reg_coeff[44]), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_n111) );
  INV_X1 my_filter_adder_mult_6_multiplication_mult_21_U217 ( .A(
        my_filter_q_reg_coeff[45]), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_n110) );
  INV_X1 my_filter_adder_mult_6_multiplication_mult_21_U216 ( .A(
        my_filter_q_reg_coeff[46]), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_n109) );
  INV_X1 my_filter_adder_mult_6_multiplication_mult_21_U215 ( .A(
        my_filter_q_reg_chain_7__8_), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_n91) );
  INV_X1 my_filter_adder_mult_6_multiplication_mult_21_U214 ( .A(
        my_filter_q_reg_chain_7__7_), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_n92) );
  INV_X1 my_filter_adder_mult_6_multiplication_mult_21_U213 ( .A(
        my_filter_q_reg_chain_7__6_), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_n93) );
  INV_X1 my_filter_adder_mult_6_multiplication_mult_21_U212 ( .A(
        my_filter_q_reg_chain_7__5_), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_n94) );
  INV_X1 my_filter_adder_mult_6_multiplication_mult_21_U211 ( .A(
        my_filter_q_reg_chain_7__4_), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_n95) );
  INV_X1 my_filter_adder_mult_6_multiplication_mult_21_U210 ( .A(
        my_filter_q_reg_chain_7__2_), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_n97) );
  INV_X1 my_filter_adder_mult_6_multiplication_mult_21_U209 ( .A(
        my_filter_q_reg_chain_7__3_), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_n96) );
  AND2_X1 my_filter_adder_mult_6_multiplication_mult_21_U208 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_13__12_), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_13__13_), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_n3) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U207 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n100), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_13__13_) );
  AND2_X1 my_filter_adder_mult_6_multiplication_mult_21_U206 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_13__11_), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_13__12_), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_n52) );
  AND2_X1 my_filter_adder_mult_6_multiplication_mult_21_U205 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_13__9_), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_13__10_), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_n50) );
  AND2_X1 my_filter_adder_mult_6_multiplication_mult_21_U204 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_13__10_), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_13__11_), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_n48) );
  AND2_X1 my_filter_adder_mult_6_multiplication_mult_21_U203 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_13__8_), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_13__9_), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_n40) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U202 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_12__11_) );
  AND2_X1 my_filter_adder_mult_6_multiplication_mult_21_U201 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_13__7_), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_13__8_), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_n46) );
  AND2_X1 my_filter_adder_mult_6_multiplication_mult_21_U200 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_13__5_), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_13__6_), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_n45) );
  AND2_X1 my_filter_adder_mult_6_multiplication_mult_21_U199 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_13__3_), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_13__4_), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_n38) );
  AND2_X1 my_filter_adder_mult_6_multiplication_mult_21_U198 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_13__1_), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_13__2_), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_n44) );
  AND2_X1 my_filter_adder_mult_6_multiplication_mult_21_U197 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_13__6_), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_13__7_), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_n39) );
  AND2_X1 my_filter_adder_mult_6_multiplication_mult_21_U196 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_13__4_), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_13__5_), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_n37) );
  AND2_X1 my_filter_adder_mult_6_multiplication_mult_21_U195 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_13__2_), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_13__3_), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_n36) );
  AND2_X1 my_filter_adder_mult_6_multiplication_mult_21_U194 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_13__0_), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_13__1_), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_n35) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U193 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_12__1_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U192 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_10__0_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U191 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_11__0_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U190 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_11__1_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U189 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_10__1_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U188 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_8__0_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U187 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n113), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_9__0_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U186 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n112), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_9__1_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U185 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n110), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_9__3_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U184 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_8__1_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U183 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_8__3_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U182 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_6__0_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U181 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_7__0_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U180 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_7__1_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U179 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_7__3_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U178 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_7__4_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U177 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_7__5_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U176 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_6__1_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U175 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_6__3_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U174 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_6__5_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U173 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_4__0_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U172 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_5__0_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U171 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_5__1_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U170 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_5__3_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U169 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_5__4_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U168 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_5__5_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U167 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_5__6_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U166 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_4__1_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U165 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_4__3_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U164 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_4__5_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U163 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_2__0_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U162 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_3__0_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U161 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_3__1_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U160 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_3__3_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U159 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_3__4_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U158 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_3__5_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U157 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_3__6_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U156 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_3__7_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U155 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_12__9_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U154 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_12__10_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U153 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_11__10_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U152 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_11__11_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U151 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_12__7_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U150 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_12__8_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U149 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_10__11_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U148 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_11__8_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U147 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_11__9_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U146 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_12__5_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U145 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_12__6_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U144 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_10__9_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U143 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_10__10_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U142 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_11__6_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U141 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_11__7_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U140 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n103), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_9__10_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U139 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n102), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_9__11_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U138 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_12__2_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U137 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_12__3_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U136 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_12__4_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U135 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_10__7_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U134 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_10__8_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U133 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_8__11_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U132 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_11__3_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U131 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_11__4_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U130 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_11__5_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U129 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n105), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_9__8_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U128 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n104), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_9__9_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U127 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_10__4_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U126 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_10__5_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U125 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_10__6_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U124 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_8__9_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U123 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_8__10_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U122 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_11__2_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U121 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n108), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_9__5_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U120 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n107), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_9__6_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U119 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n106), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_9__7_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U118 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_7__10_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U117 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_7__11_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U116 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_10__2_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U115 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_10__3_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U114 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_8__6_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U113 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_8__7_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U112 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_8__8_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U111 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_6__11_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U110 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n111), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_9__2_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U109 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n109), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_9__4_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U108 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_7__7_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U107 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_7__8_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U106 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_7__9_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U105 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_8__2_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U104 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_8__4_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U103 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_8__5_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U102 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_6__8_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U101 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_6__9_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U100 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_6__10_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U99 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_7__2_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U98 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_7__6_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U97 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_5__9_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U96 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_5__10_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U95 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_5__11_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U94 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_6__2_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U93 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_6__4_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U92 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_6__6_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U91 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_6__7_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U90 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_4__10_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U89 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_4__11_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U88 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_5__2_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U87 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_5__7_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U86 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_5__8_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U85 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_3__11_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U84 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_4__2_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U83 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_4__4_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U82 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_4__6_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U81 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_4__7_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U80 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_4__8_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U79 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_4__9_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U78 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_3__2_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U77 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_3__8_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U76 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_3__9_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U75 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_3__10_) );
  AND2_X1 my_filter_adder_mult_6_multiplication_mult_21_U74 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_ab_0__2_), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_ab_1__1_), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_n14) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U73 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_2__1_) );
  AND2_X1 my_filter_adder_mult_6_multiplication_mult_21_U72 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_ab_0__3_), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_ab_1__2_), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_n13) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U71 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_2__2_) );
  AND2_X1 my_filter_adder_mult_6_multiplication_mult_21_U70 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_ab_0__4_), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_ab_1__3_), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_n12) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U69 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_2__3_) );
  AND2_X1 my_filter_adder_mult_6_multiplication_mult_21_U68 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_ab_0__5_), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_ab_1__4_), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_n11) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U67 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_2__4_) );
  AND2_X1 my_filter_adder_mult_6_multiplication_mult_21_U66 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_ab_0__6_), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_ab_1__5_), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_n10) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U65 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_2__5_) );
  AND2_X1 my_filter_adder_mult_6_multiplication_mult_21_U64 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_ab_0__7_), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_ab_1__6_), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_n9) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U63 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_2__6_) );
  AND2_X1 my_filter_adder_mult_6_multiplication_mult_21_U62 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_ab_0__8_), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_ab_1__7_), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_n8) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U61 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_2__7_) );
  AND2_X1 my_filter_adder_mult_6_multiplication_mult_21_U60 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_ab_0__9_), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_ab_1__8_), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_n7) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U59 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_2__8_) );
  AND2_X1 my_filter_adder_mult_6_multiplication_mult_21_U58 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_ab_0__10_), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_ab_1__9_), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_n6) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U57 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_2__9_) );
  AND2_X1 my_filter_adder_mult_6_multiplication_mult_21_U56 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_ab_0__11_), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_ab_1__10_), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_n5) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U55 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_2__10_) );
  AND2_X1 my_filter_adder_mult_6_multiplication_mult_21_U54 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_ab_0__12_), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_ab_1__11_), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_n4) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U52 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_2__11_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U50 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_1__12_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U48 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_1__2_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U46 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_1__3_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U45 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_1__4_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U44 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_1__5_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U40 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_1__6_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U39 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_1__7_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U38 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_1__8_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U37 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_1__9_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U36 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_1__10_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U35 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_1__11_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U14 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_0__2_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U13 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_0__3_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U12 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_0__4_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U11 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_0__5_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U10 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_0__6_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U9 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_0__7_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U8 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_0__8_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U7 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_0__9_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U6 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_0__10_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U5 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_0__11_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U4 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_0__12_) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U3 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n98), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n112), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_ab_1__1_) );
  INV_X1 my_filter_adder_mult_6_multiplication_mult_21_U2 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_13__13_), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_n85) );
  XOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U51 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_13__12_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_13__13_), .Z(
        my_filter_adder_mult_6_multiplication_mult_21_n51) );
  XOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U49 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_13__10_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_13__11_), .Z(
        my_filter_adder_mult_6_multiplication_mult_21_n49) );
  XOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U47 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_13__11_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_13__12_), .Z(
        my_filter_adder_mult_6_multiplication_mult_21_n47) );
  XOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U43 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_13__5_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_13__6_), .Z(
        my_filter_adder_mult_6_multiplication_mult_21_n43) );
  XOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U42 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_13__3_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_13__4_), .Z(
        my_filter_adder_mult_6_multiplication_mult_21_n42) );
  XOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U41 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_13__1_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_13__2_), .Z(
        my_filter_adder_mult_6_multiplication_mult_21_n41) );
  XOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U34 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_13__8_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_13__9_), .Z(
        my_filter_adder_mult_6_multiplication_mult_21_n34) );
  XOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U33 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_13__9_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_13__10_), .Z(
        my_filter_adder_mult_6_multiplication_mult_21_n33) );
  XOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U32 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_13__6_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_13__7_), .Z(
        my_filter_adder_mult_6_multiplication_mult_21_n32) );
  XOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U31 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_13__7_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_13__8_), .Z(
        my_filter_adder_mult_6_multiplication_mult_21_n31) );
  XOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U30 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_13__4_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_13__5_), .Z(
        my_filter_adder_mult_6_multiplication_mult_21_n30) );
  XOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U29 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_13__2_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_13__3_), .Z(
        my_filter_adder_mult_6_multiplication_mult_21_n29) );
  XOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U28 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_13__0_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_13__1_), .Z(
        my_filter_adder_mult_6_multiplication_mult_21_n28) );
  XOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U26 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_1__1_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_ab_0__2_), .Z(
        my_filter_adder_mult_6_multiplication_mult_21_n27) );
  XOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U25 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_1__12_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_ab_0__13_), .Z(
        my_filter_adder_mult_6_multiplication_mult_21_n26) );
  XOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U24 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_1__2_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_ab_0__3_), .Z(
        my_filter_adder_mult_6_multiplication_mult_21_n25) );
  XOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U23 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_1__3_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_ab_0__4_), .Z(
        my_filter_adder_mult_6_multiplication_mult_21_n24) );
  XOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U22 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_1__4_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_ab_0__5_), .Z(
        my_filter_adder_mult_6_multiplication_mult_21_n23) );
  XOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U21 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_1__5_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_ab_0__6_), .Z(
        my_filter_adder_mult_6_multiplication_mult_21_n22) );
  XOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U20 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_1__6_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_ab_0__7_), .Z(
        my_filter_adder_mult_6_multiplication_mult_21_n21) );
  XOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U19 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_1__7_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_ab_0__8_), .Z(
        my_filter_adder_mult_6_multiplication_mult_21_n20) );
  XOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U18 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_1__8_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_ab_0__9_), .Z(
        my_filter_adder_mult_6_multiplication_mult_21_n19) );
  XOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U17 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_1__9_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_ab_0__10_), .Z(
        my_filter_adder_mult_6_multiplication_mult_21_n18) );
  XOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U16 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_1__10_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_ab_0__11_), .Z(
        my_filter_adder_mult_6_multiplication_mult_21_n17) );
  XOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_U15 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_1__11_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_ab_0__12_), .Z(
        my_filter_adder_mult_6_multiplication_mult_21_n16) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S3_2_12 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_2__12_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_n15), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_ab_1__13_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_2__12_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_2__12_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_2_11 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_2__11_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_n4), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_n26), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_2__11_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_2__11_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_2_10 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_2__10_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_n5), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_n16), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_2__10_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_2__10_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_2_9 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_2__9_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_n6), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_n17), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_2__9_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_2__9_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_2_8 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_2__8_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_n7), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_n18), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_2__8_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_2__8_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_2_7 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_2__7_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_n8), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_n19), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_2__7_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_2__7_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_2_6 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_2__6_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_n9), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_n20), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_2__6_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_2__6_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_2_5 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_2__5_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_n10), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_n21), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_2__5_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_2__5_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_2_4 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_2__4_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_n11), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_n22), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_2__4_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_2__4_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_2_3 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_2__3_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_n12), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_n23), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_2__3_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_2__3_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_2_2 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_2__2_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_n13), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_n24), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_2__2_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_2__2_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_2_1 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_2__1_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_n14), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_n25), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_2__1_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_2__1_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S1_2_0 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_2__0_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_1__0_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_n27), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_2__0_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_A1_0_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S3_3_12 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_3__12_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_2__12_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_ab_2__13_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_3__12_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_3__12_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_3_11 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_3__11_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_2__11_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_2__12_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_3__11_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_3__11_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_3_10 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_3__10_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_2__10_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_2__11_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_3__10_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_3__10_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_3_9 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_3__9_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_2__9_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_2__10_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_3__9_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_3__9_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_3_8 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_3__8_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_2__8_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_2__9_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_3__8_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_3__8_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_3_7 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_3__7_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_2__7_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_2__8_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_3__7_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_3__7_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_3_6 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_3__6_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_2__6_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_2__7_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_3__6_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_3__6_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_3_5 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_3__5_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_2__5_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_2__6_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_3__5_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_3__5_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_3_4 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_3__4_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_2__4_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_2__5_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_3__4_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_3__4_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_3_3 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_3__3_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_2__3_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_2__4_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_3__3_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_3__3_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_3_2 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_3__2_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_2__2_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_2__3_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_3__2_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_3__2_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_3_1 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_3__1_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_2__1_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_2__2_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_3__1_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_3__1_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S1_3_0 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_3__0_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_2__0_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_2__1_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_3__0_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_A1_1_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S3_4_12 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_4__12_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_3__12_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_ab_3__13_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_4__12_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_4__12_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_4_11 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_4__11_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_3__11_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_3__12_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_4__11_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_4__11_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_4_10 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_4__10_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_3__10_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_3__11_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_4__10_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_4__10_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_4_9 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_4__9_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_3__9_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_3__10_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_4__9_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_4__9_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_4_8 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_4__8_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_3__8_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_3__9_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_4__8_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_4__8_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_4_7 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_4__7_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_3__7_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_3__8_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_4__7_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_4__7_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_4_6 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_4__6_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_3__6_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_3__7_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_4__6_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_4__6_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_4_5 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_4__5_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_3__5_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_3__6_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_4__5_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_4__5_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_4_4 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_4__4_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_3__4_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_3__5_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_4__4_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_4__4_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_4_3 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_4__3_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_3__3_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_3__4_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_4__3_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_4__3_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_4_2 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_4__2_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_3__2_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_3__3_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_4__2_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_4__2_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_4_1 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_4__1_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_3__1_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_3__2_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_4__1_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_4__1_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S1_4_0 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_4__0_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_3__0_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_3__1_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_4__0_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_A1_2_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S3_5_12 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_5__12_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_4__12_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_ab_4__13_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_5__12_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_5__12_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_5_11 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_5__11_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_4__11_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_4__12_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_5__11_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_5__11_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_5_10 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_5__10_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_4__10_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_4__11_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_5__10_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_5__10_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_5_9 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_5__9_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_4__9_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_4__10_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_5__9_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_5__9_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_5_8 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_5__8_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_4__8_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_4__9_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_5__8_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_5__8_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_5_7 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_5__7_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_4__7_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_4__8_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_5__7_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_5__7_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_5_6 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_5__6_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_4__6_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_4__7_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_5__6_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_5__6_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_5_5 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_5__5_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_4__5_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_4__6_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_5__5_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_5__5_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_5_4 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_5__4_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_4__4_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_4__5_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_5__4_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_5__4_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_5_3 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_5__3_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_4__3_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_4__4_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_5__3_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_5__3_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_5_2 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_5__2_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_4__2_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_4__3_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_5__2_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_5__2_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_5_1 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_5__1_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_4__1_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_4__2_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_5__1_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_5__1_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S1_5_0 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_5__0_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_4__0_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_4__1_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_5__0_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_A1_3_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S3_6_12 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_6__12_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_5__12_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_ab_5__13_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_6__12_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_6__12_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_6_11 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_6__11_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_5__11_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_5__12_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_6__11_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_6__11_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_6_10 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_6__10_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_5__10_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_5__11_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_6__10_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_6__10_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_6_9 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_6__9_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_5__9_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_5__10_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_6__9_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_6__9_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_6_8 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_6__8_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_5__8_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_5__9_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_6__8_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_6__8_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_6_7 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_6__7_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_5__7_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_5__8_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_6__7_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_6__7_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_6_6 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_6__6_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_5__6_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_5__7_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_6__6_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_6__6_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_6_5 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_6__5_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_5__5_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_5__6_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_6__5_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_6__5_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_6_4 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_6__4_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_5__4_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_5__5_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_6__4_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_6__4_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_6_3 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_6__3_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_5__3_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_5__4_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_6__3_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_6__3_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_6_2 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_6__2_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_5__2_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_5__3_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_6__2_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_6__2_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_6_1 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_6__1_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_5__1_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_5__2_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_6__1_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_6__1_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S1_6_0 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_6__0_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_5__0_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_5__1_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_6__0_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_A1_4_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S3_7_12 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_7__12_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_6__12_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_ab_6__13_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_7__12_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_7__12_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_7_11 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_7__11_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_6__11_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_6__12_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_7__11_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_7__11_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_7_10 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_7__10_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_6__10_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_6__11_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_7__10_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_7__10_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_7_9 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_7__9_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_6__9_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_6__10_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_7__9_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_7__9_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_7_8 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_7__8_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_6__8_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_6__9_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_7__8_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_7__8_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_7_7 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_7__7_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_6__7_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_6__8_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_7__7_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_7__7_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_7_6 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_7__6_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_6__6_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_6__7_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_7__6_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_7__6_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_7_5 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_7__5_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_6__5_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_6__6_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_7__5_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_7__5_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_7_4 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_7__4_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_6__4_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_6__5_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_7__4_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_7__4_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_7_3 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_7__3_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_6__3_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_6__4_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_7__3_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_7__3_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_7_2 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_7__2_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_6__2_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_6__3_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_7__2_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_7__2_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_7_1 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_7__1_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_6__1_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_6__2_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_7__1_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_7__1_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S1_7_0 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_7__0_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_6__0_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_6__1_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_7__0_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_A1_5_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S3_8_12 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_8__12_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_7__12_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_ab_7__13_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_8__12_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_8__12_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_8_11 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_8__11_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_7__11_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_7__12_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_8__11_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_8__11_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_8_10 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_8__10_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_7__10_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_7__11_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_8__10_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_8__10_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_8_9 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_8__9_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_7__9_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_7__10_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_8__9_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_8__9_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_8_8 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_8__8_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_7__8_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_7__9_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_8__8_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_8__8_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_8_7 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_8__7_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_7__7_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_7__8_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_8__7_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_8__7_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_8_6 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_8__6_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_7__6_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_7__7_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_8__6_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_8__6_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_8_5 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_8__5_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_7__5_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_7__6_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_8__5_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_8__5_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_8_4 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_8__4_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_7__4_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_7__5_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_8__4_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_8__4_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_8_3 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_8__3_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_7__3_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_7__4_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_8__3_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_8__3_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_8_2 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_8__2_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_7__2_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_7__3_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_8__2_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_8__2_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_8_1 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_8__1_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_7__1_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_7__2_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_8__1_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_8__1_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S1_8_0 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_8__0_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_7__0_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_7__1_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_8__0_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_A1_6_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S3_9_12 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_9__12_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_8__12_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_ab_8__13_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_9__12_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_9__12_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_9_11 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_9__11_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_8__11_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_8__12_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_9__11_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_9__11_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_9_10 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_9__10_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_8__10_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_8__11_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_9__10_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_9__10_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_9_9 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_9__9_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_8__9_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_8__10_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_9__9_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_9__9_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_9_8 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_9__8_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_8__8_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_8__9_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_9__8_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_9__8_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_9_7 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_9__7_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_8__7_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_8__8_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_9__7_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_9__7_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_9_6 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_9__6_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_8__6_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_8__7_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_9__6_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_9__6_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_9_5 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_9__5_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_8__5_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_8__6_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_9__5_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_9__5_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_9_4 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_9__4_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_8__4_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_8__5_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_9__4_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_9__4_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_9_3 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_9__3_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_8__3_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_8__4_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_9__3_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_9__3_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_9_2 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_9__2_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_8__2_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_8__3_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_9__2_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_9__2_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_9_1 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_9__1_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_8__1_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_8__2_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_9__1_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_9__1_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S1_9_0 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_9__0_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_8__0_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_8__1_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_9__0_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_A1_7_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S3_10_12 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_10__12_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_9__12_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_ab_9__13_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_10__12_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_10__12_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_10_11 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_10__11_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_9__11_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_9__12_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_10__11_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_10__11_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_10_10 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_10__10_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_9__10_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_9__11_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_10__10_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_10__10_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_10_9 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_10__9_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_9__9_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_9__10_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_10__9_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_10__9_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_10_8 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_10__8_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_9__8_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_9__9_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_10__8_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_10__8_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_10_7 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_10__7_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_9__7_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_9__8_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_10__7_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_10__7_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_10_6 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_10__6_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_9__6_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_9__7_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_10__6_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_10__6_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_10_5 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_10__5_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_9__5_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_9__6_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_10__5_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_10__5_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_10_4 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_10__4_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_9__4_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_9__5_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_10__4_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_10__4_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_10_3 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_10__3_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_9__3_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_9__4_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_10__3_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_10__3_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_10_2 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_10__2_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_9__2_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_9__3_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_10__2_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_10__2_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_10_1 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_10__1_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_9__1_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_9__2_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_10__1_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_10__1_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S1_10_0 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_10__0_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_9__0_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_9__1_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_10__0_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_A1_8_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S3_11_12 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_11__12_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_10__12_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_ab_10__13_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_11__12_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_11__12_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_11_11 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_11__11_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_10__11_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_10__12_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_11__11_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_11__11_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_11_10 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_11__10_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_10__10_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_10__11_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_11__10_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_11__10_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_11_9 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_11__9_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_10__9_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_10__10_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_11__9_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_11__9_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_11_8 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_11__8_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_10__8_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_10__9_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_11__8_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_11__8_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_11_7 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_11__7_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_10__7_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_10__8_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_11__7_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_11__7_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_11_6 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_11__6_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_10__6_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_10__7_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_11__6_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_11__6_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_11_5 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_11__5_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_10__5_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_10__6_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_11__5_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_11__5_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_11_4 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_11__4_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_10__4_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_10__5_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_11__4_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_11__4_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_11_3 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_11__3_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_10__3_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_10__4_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_11__3_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_11__3_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_11_2 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_11__2_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_10__2_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_10__3_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_11__2_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_11__2_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_11_1 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_11__1_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_10__1_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_10__2_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_11__1_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_11__1_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S1_11_0 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_11__0_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_10__0_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_10__1_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_11__0_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_A1_9_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S3_12_12 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_12__12_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_11__12_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_ab_11__13_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_12__12_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_12__12_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_12_11 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_12__11_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_11__11_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_11__12_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_12__11_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_12__11_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_12_10 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_12__10_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_11__10_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_11__11_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_12__10_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_12__10_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_12_9 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_12__9_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_11__9_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_11__10_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_12__9_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_12__9_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_12_8 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_12__8_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_11__8_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_11__9_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_12__8_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_12__8_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_12_7 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_12__7_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_11__7_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_11__8_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_12__7_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_12__7_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_12_6 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_12__6_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_11__6_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_11__7_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_12__6_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_12__6_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_12_5 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_12__5_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_11__5_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_11__6_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_12__5_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_12__5_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_12_4 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_12__4_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_11__4_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_11__5_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_12__4_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_12__4_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_12_3 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_12__3_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_11__3_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_11__4_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_12__3_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_12__3_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_12_2 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_12__2_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_11__2_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_11__3_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_12__2_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_12__2_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S2_12_1 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_12__1_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_11__1_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_11__2_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_12__1_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_12__1_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S1_12_0 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_12__0_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_11__0_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_11__1_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_12__0_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_A1_10_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S14_13 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_n86), .B(
        my_filter_adder_mult_6_multiplication_mult_21_n100), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_ab_13__13_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_13__13_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_13__13_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S5_12 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_13__12_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_12__12_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_ab_12__13_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_13__12_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_13__12_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S4_11 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_13__11_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_12__11_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_12__12_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_13__11_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_13__11_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S4_10 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_13__10_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_12__10_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_12__11_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_13__10_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_13__10_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S4_9 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_13__9_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_12__9_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_12__10_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_13__9_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_13__9_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S4_8 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_13__8_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_12__8_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_12__9_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_13__8_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_13__8_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S4_7 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_13__7_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_12__7_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_12__8_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_13__7_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_13__7_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S4_6 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_13__6_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_12__6_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_12__7_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_13__6_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_13__6_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S4_5 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_13__5_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_12__5_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_12__6_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_13__5_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_13__5_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S4_4 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_13__4_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_12__4_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_12__5_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_13__4_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_13__4_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S4_3 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_13__3_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_12__3_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_12__4_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_13__3_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_13__3_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S4_2 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_13__2_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_12__2_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_12__3_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_13__2_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_13__2_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S4_1 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_13__1_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_12__1_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_12__2_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_13__1_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_13__1_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S4_0 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_ab_13__0_), .B(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_12__0_), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_12__1_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_CARRYB_13__0_), .S(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_13__0_) );
  FA_X1 my_filter_adder_mult_6_multiplication_mult_21_S14_13_0 ( .A(
        my_filter_q_reg_chain_7__13_), .B(my_filter_q_reg_coeff[55]), .CI(
        my_filter_adder_mult_6_multiplication_mult_21_SUMB_13__0_), .CO(
        my_filter_adder_mult_6_multiplication_mult_21_A2_12_), .S(
        my_filter_adder_mult_6_res_mult[0]) );
  NAND2_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U72 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_A2_12_), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n28), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n56) );
  OAI21_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U71 ( .B1(
        my_filter_adder_mult_6_multiplication_mult_21_A2_12_), .B2(
        my_filter_adder_mult_6_multiplication_mult_21_n28), .A(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n56), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n59) );
  INV_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U70 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n59), .ZN(
        my_filter_adder_mult_6_res_mult[1]) );
  AND2_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U69 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n50), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n49), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n20) );
  NAND2_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U68 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n48), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n47), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n17) );
  NAND2_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U66 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n40), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n33), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n25) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U65 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n48), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n47), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n15) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U64 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n40), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n33), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n23) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U63 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n50), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n49), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n21) );
  AND2_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U61 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n46), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n34), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n28) );
  AND2_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U60 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n45), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n32), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n36) );
  AND2_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U59 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n38), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n30), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n44) );
  AND2_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U58 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n44), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n29), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n52) );
  NAND2_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U56 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n39), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n31), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n33) );
  NAND2_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U55 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n37), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n43), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n41) );
  NAND2_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U54 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n36), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n42), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n49) );
  NAND2_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U53 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n35), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n41), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n57) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U51 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n39), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n31), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n31) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U50 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n37), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n43), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n39) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U49 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n36), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n42), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n47) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U48 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n35), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n41), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n55) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U46 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n46), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n34), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n29) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U45 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n45), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n32), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n37) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U44 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n38), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n30), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n45) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U43 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_n44), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_n29), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n53) );
  OAI21_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U41 ( .B1(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n55), .B2(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n56), .A(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n57), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n51) );
  INV_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U40 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n55), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n60) );
  NAND2_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U39 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n60), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n57), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n58) );
  OAI21_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U38 ( .B1(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n15), .B2(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n16), .A(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n17), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n13) );
  OAI21_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U36 ( .B1(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n23), .B2(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n24), .A(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n25), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n19) );
  OAI21_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U35 ( .B1(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n31), .B2(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n32), .A(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n33), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n27) );
  OAI21_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U34 ( .B1(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n39), .B2(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n40), .A(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n41), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n35) );
  OAI21_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U33 ( .B1(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n47), .B2(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n48), .A(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n49), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n43) );
  INV_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U31 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n21), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n63) );
  AOI21_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U30 ( .B1(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n63), .B2(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n19), .A(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n20), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n16) );
  INV_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U29 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n29), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n71) );
  AOI21_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U28 ( .B1(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n71), .B2(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n27), .A(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n28), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n24) );
  INV_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U26 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n37), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n69) );
  AOI21_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U25 ( .B1(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n69), .B2(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n35), .A(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n36), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n32) );
  INV_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U24 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n45), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n67) );
  AOI21_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U23 ( .B1(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n67), .B2(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n43), .A(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n44), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n40) );
  INV_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U21 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n53), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n65) );
  AOI21_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U20 ( .B1(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n65), .B2(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n51), .A(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n52), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n48) );
  INV_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U19 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n15), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n62) );
  NAND2_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U18 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n62), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n17), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n18) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U16 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n20), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n21), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n22) );
  INV_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U13 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n23), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n64) );
  NAND2_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U12 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n64), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n25), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n26) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U11 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n28), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n29), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n30) );
  INV_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U10 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n31), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n70) );
  NAND2_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U9 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n70), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n33), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n34) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U8 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n36), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n37), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n38) );
  INV_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U7 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n39), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n68) );
  NAND2_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U6 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n68), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n41), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n42) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U5 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n44), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n45), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n46) );
  INV_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U4 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n47), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n66) );
  NAND2_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U3 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n66), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n49), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n50) );
  NOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U2 ( .A1(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n52), .A2(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n53), .ZN(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n54) );
  XOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U67 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n56), .B(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n58), .Z(
        my_filter_adder_mult_6_res_mult[2]) );
  XOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U62 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n51), .B(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n54), .Z(
        my_filter_adder_mult_6_res_mult[3]) );
  XOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U57 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n50), .B(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n48), .Z(
        my_filter_adder_mult_6_res_mult[4]) );
  XOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U52 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n43), .B(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n46), .Z(
        my_filter_adder_mult_6_res_mult[5]) );
  XOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U47 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n42), .B(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n40), .Z(
        my_filter_adder_mult_6_res_mult[6]) );
  XOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U42 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n35), .B(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n38), .Z(
        my_filter_adder_mult_6_res_mult[7]) );
  XOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U37 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n34), .B(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n32), .Z(
        my_filter_adder_mult_6_res_mult[8]) );
  XOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U32 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n27), .B(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n30), .Z(
        my_filter_adder_mult_6_res_mult[9]) );
  XOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U27 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n26), .B(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n24), .Z(
        my_filter_adder_mult_6_res_mult[10]) );
  XOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U22 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n19), .B(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n22), .Z(
        my_filter_adder_mult_6_res_mult[11]) );
  XOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U17 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n18), .B(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n16), .Z(
        my_filter_adder_mult_6_res_mult[12]) );
  XOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U15 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_n52), .B(
        my_filter_adder_mult_6_multiplication_mult_21_n51), .Z(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n14) );
  XOR2_X1 my_filter_adder_mult_6_multiplication_mult_21_FS_1_U14 ( .A(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n13), .B(
        my_filter_adder_mult_6_multiplication_mult_21_FS_1_n14), .Z(
        my_filter_adder_mult_6_res_mult[13]) );
  AND2_X1 my_filter_adder_mult_6_addition_add_19_U1 ( .A1(
        my_filter_data_sum[56]), .A2(my_filter_adder_mult_6_res_mult[0]), .ZN(
        my_filter_adder_mult_6_addition_add_19_n1) );
  XOR2_X1 my_filter_adder_mult_6_addition_add_19_U2 ( .A(
        my_filter_data_sum[56]), .B(my_filter_adder_mult_6_res_mult[0]), .Z(
        my_filter_data_sum[42]) );
  FA_X1 my_filter_adder_mult_6_addition_add_19_U1_1 ( .A(
        my_filter_adder_mult_6_res_mult[1]), .B(my_filter_data_sum[57]), .CI(
        my_filter_adder_mult_6_addition_add_19_n1), .CO(
        my_filter_adder_mult_6_addition_add_19_carry[2]), .S(
        my_filter_data_sum[43]) );
  FA_X1 my_filter_adder_mult_6_addition_add_19_U1_2 ( .A(
        my_filter_adder_mult_6_res_mult[2]), .B(my_filter_data_sum[58]), .CI(
        my_filter_adder_mult_6_addition_add_19_carry[2]), .CO(
        my_filter_adder_mult_6_addition_add_19_carry[3]), .S(
        my_filter_data_sum[44]) );
  FA_X1 my_filter_adder_mult_6_addition_add_19_U1_3 ( .A(
        my_filter_adder_mult_6_res_mult[3]), .B(my_filter_data_sum[59]), .CI(
        my_filter_adder_mult_6_addition_add_19_carry[3]), .CO(
        my_filter_adder_mult_6_addition_add_19_carry[4]), .S(
        my_filter_data_sum[45]) );
  FA_X1 my_filter_adder_mult_6_addition_add_19_U1_4 ( .A(
        my_filter_adder_mult_6_res_mult[4]), .B(my_filter_data_sum[60]), .CI(
        my_filter_adder_mult_6_addition_add_19_carry[4]), .CO(
        my_filter_adder_mult_6_addition_add_19_carry[5]), .S(
        my_filter_data_sum[46]) );
  FA_X1 my_filter_adder_mult_6_addition_add_19_U1_5 ( .A(
        my_filter_adder_mult_6_res_mult[5]), .B(my_filter_data_sum[61]), .CI(
        my_filter_adder_mult_6_addition_add_19_carry[5]), .CO(
        my_filter_adder_mult_6_addition_add_19_carry[6]), .S(
        my_filter_data_sum[47]) );
  FA_X1 my_filter_adder_mult_6_addition_add_19_U1_6 ( .A(
        my_filter_adder_mult_6_res_mult[6]), .B(my_filter_data_sum[62]), .CI(
        my_filter_adder_mult_6_addition_add_19_carry[6]), .CO(
        my_filter_adder_mult_6_addition_add_19_carry[7]), .S(
        my_filter_data_sum[48]) );
  FA_X1 my_filter_adder_mult_6_addition_add_19_U1_7 ( .A(
        my_filter_adder_mult_6_res_mult[7]), .B(my_filter_data_sum[63]), .CI(
        my_filter_adder_mult_6_addition_add_19_carry[7]), .CO(
        my_filter_adder_mult_6_addition_add_19_carry[8]), .S(
        my_filter_data_sum[49]) );
  FA_X1 my_filter_adder_mult_6_addition_add_19_U1_8 ( .A(
        my_filter_adder_mult_6_res_mult[8]), .B(my_filter_data_sum[64]), .CI(
        my_filter_adder_mult_6_addition_add_19_carry[8]), .CO(
        my_filter_adder_mult_6_addition_add_19_carry[9]), .S(
        my_filter_data_sum[50]) );
  FA_X1 my_filter_adder_mult_6_addition_add_19_U1_9 ( .A(
        my_filter_adder_mult_6_res_mult[9]), .B(my_filter_data_sum[65]), .CI(
        my_filter_adder_mult_6_addition_add_19_carry[9]), .CO(
        my_filter_adder_mult_6_addition_add_19_carry[10]), .S(
        my_filter_data_sum[51]) );
  FA_X1 my_filter_adder_mult_6_addition_add_19_U1_10 ( .A(
        my_filter_adder_mult_6_res_mult[10]), .B(my_filter_data_sum[66]), .CI(
        my_filter_adder_mult_6_addition_add_19_carry[10]), .CO(
        my_filter_adder_mult_6_addition_add_19_carry[11]), .S(
        my_filter_data_sum[52]) );
  FA_X1 my_filter_adder_mult_6_addition_add_19_U1_11 ( .A(
        my_filter_adder_mult_6_res_mult[11]), .B(my_filter_data_sum[67]), .CI(
        my_filter_adder_mult_6_addition_add_19_carry[11]), .CO(
        my_filter_adder_mult_6_addition_add_19_carry[12]), .S(
        my_filter_data_sum[53]) );
  FA_X1 my_filter_adder_mult_6_addition_add_19_U1_12 ( .A(
        my_filter_adder_mult_6_res_mult[12]), .B(my_filter_data_sum[68]), .CI(
        my_filter_adder_mult_6_addition_add_19_carry[12]), .CO(
        my_filter_adder_mult_6_addition_add_19_carry[13]), .S(
        my_filter_data_sum[54]) );
  FA_X1 my_filter_adder_mult_6_addition_add_19_U1_13 ( .A(
        my_filter_adder_mult_6_res_mult[13]), .B(my_filter_data_sum[69]), .CI(
        my_filter_adder_mult_6_addition_add_19_carry[13]), .S(
        my_filter_data_sum[55]) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U276 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_12__12_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U275 ( .A1(
        my_filter_q_reg_chain_8__11_), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_11__13_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U274 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_11__12_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U273 ( .A1(
        my_filter_q_reg_chain_8__10_), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_10__13_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U272 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_10__12_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U271 ( .A1(
        my_filter_q_reg_chain_8__9_), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_9__13_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U270 ( .A1(
        my_filter_q_reg_coeff[39]), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_13__11_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U269 ( .A1(
        my_filter_q_reg_coeff[38]), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_13__10_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U268 ( .A1(
        my_filter_q_reg_coeff[37]), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_13__9_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U267 ( .A1(
        my_filter_q_reg_coeff[40]), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_13__12_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U266 ( .A1(
        my_filter_q_reg_chain_8__12_), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_12__13_) );
  INV_X1 my_filter_adder_mult_7_multiplication_mult_21_U265 ( .A(
        my_filter_q_reg_chain_8__9_), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_n90) );
  INV_X1 my_filter_adder_mult_7_multiplication_mult_21_U264 ( .A(
        my_filter_q_reg_chain_8__12_), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_n87) );
  INV_X1 my_filter_adder_mult_7_multiplication_mult_21_U263 ( .A(
        my_filter_q_reg_chain_8__11_), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_n88) );
  INV_X1 my_filter_adder_mult_7_multiplication_mult_21_U262 ( .A(
        my_filter_q_reg_chain_8__10_), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_n89) );
  INV_X1 my_filter_adder_mult_7_multiplication_mult_21_U261 ( .A(
        my_filter_q_reg_chain_8__8_), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_n91) );
  INV_X1 my_filter_adder_mult_7_multiplication_mult_21_U260 ( .A(
        my_filter_q_reg_chain_8__13_), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_n86) );
  AND2_X1 my_filter_adder_mult_7_multiplication_mult_21_U259 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_ab_0__13_), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_ab_1__12_), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_n15) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U258 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_2__12_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U257 ( .A1(
        my_filter_q_reg_chain_8__1_), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_1__13_) );
  AND3_X1 my_filter_adder_mult_7_multiplication_mult_21_U256 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_ab_1__1_), .A2(
        my_filter_q_reg_coeff[28]), .A3(my_filter_q_reg_chain_8__0_), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_1__0_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U255 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_12__0_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U254 ( .A1(
        my_filter_q_reg_coeff[28]), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_13__0_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U253 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n101), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_9__12_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U252 ( .A1(
        my_filter_q_reg_chain_8__8_), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_8__13_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U251 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_8__12_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U250 ( .A1(
        my_filter_q_reg_chain_8__7_), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_7__13_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U249 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_7__12_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U248 ( .A1(
        my_filter_q_reg_chain_8__6_), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_6__13_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U247 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_6__12_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U246 ( .A1(
        my_filter_q_reg_chain_8__5_), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_5__13_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U245 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_5__12_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U244 ( .A1(
        my_filter_q_reg_chain_8__4_), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_4__13_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U243 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_4__12_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U242 ( .A1(
        my_filter_q_reg_chain_8__3_), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_3__13_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U241 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_3__12_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U240 ( .A1(
        my_filter_q_reg_chain_8__2_), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_2__13_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U239 ( .A1(
        my_filter_q_reg_coeff[36]), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_13__8_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U238 ( .A1(
        my_filter_q_reg_coeff[34]), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_13__6_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U237 ( .A1(
        my_filter_q_reg_coeff[35]), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_13__7_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U236 ( .A1(
        my_filter_q_reg_coeff[32]), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_13__4_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U235 ( .A1(
        my_filter_q_reg_coeff[33]), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_13__5_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U234 ( .A1(
        my_filter_q_reg_coeff[29]), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_13__1_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U233 ( .A1(
        my_filter_q_reg_coeff[30]), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_13__2_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U232 ( .A1(
        my_filter_q_reg_coeff[31]), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_13__3_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U231 ( .A1(
        my_filter_q_reg_chain_8__0_), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_0__13_) );
  INV_X1 my_filter_adder_mult_7_multiplication_mult_21_U230 ( .A(
        my_filter_q_reg_coeff[41]), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_n100) );
  INV_X1 my_filter_adder_mult_7_multiplication_mult_21_U229 ( .A(
        my_filter_q_reg_coeff[28]), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_n113) );
  INV_X1 my_filter_adder_mult_7_multiplication_mult_21_U228 ( .A(
        my_filter_q_reg_chain_8__0_), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_n99) );
  INV_X1 my_filter_adder_mult_7_multiplication_mult_21_U227 ( .A(
        my_filter_q_reg_coeff[29]), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_n112) );
  INV_X1 my_filter_adder_mult_7_multiplication_mult_21_U226 ( .A(
        my_filter_q_reg_chain_8__1_), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_n98) );
  INV_X1 my_filter_adder_mult_7_multiplication_mult_21_U225 ( .A(
        my_filter_q_reg_coeff[40]), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_n101) );
  INV_X1 my_filter_adder_mult_7_multiplication_mult_21_U224 ( .A(
        my_filter_q_reg_coeff[38]), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_n103) );
  INV_X1 my_filter_adder_mult_7_multiplication_mult_21_U223 ( .A(
        my_filter_q_reg_coeff[39]), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_n102) );
  INV_X1 my_filter_adder_mult_7_multiplication_mult_21_U222 ( .A(
        my_filter_q_reg_coeff[36]), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_n105) );
  INV_X1 my_filter_adder_mult_7_multiplication_mult_21_U221 ( .A(
        my_filter_q_reg_coeff[37]), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_n104) );
  INV_X1 my_filter_adder_mult_7_multiplication_mult_21_U220 ( .A(
        my_filter_q_reg_coeff[33]), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_n108) );
  INV_X1 my_filter_adder_mult_7_multiplication_mult_21_U219 ( .A(
        my_filter_q_reg_coeff[34]), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_n107) );
  INV_X1 my_filter_adder_mult_7_multiplication_mult_21_U218 ( .A(
        my_filter_q_reg_coeff[35]), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_n106) );
  INV_X1 my_filter_adder_mult_7_multiplication_mult_21_U217 ( .A(
        my_filter_q_reg_coeff[30]), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_n111) );
  INV_X1 my_filter_adder_mult_7_multiplication_mult_21_U216 ( .A(
        my_filter_q_reg_coeff[31]), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_n110) );
  INV_X1 my_filter_adder_mult_7_multiplication_mult_21_U215 ( .A(
        my_filter_q_reg_coeff[32]), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_n109) );
  INV_X1 my_filter_adder_mult_7_multiplication_mult_21_U214 ( .A(
        my_filter_q_reg_chain_8__7_), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_n92) );
  INV_X1 my_filter_adder_mult_7_multiplication_mult_21_U213 ( .A(
        my_filter_q_reg_chain_8__6_), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_n93) );
  INV_X1 my_filter_adder_mult_7_multiplication_mult_21_U212 ( .A(
        my_filter_q_reg_chain_8__5_), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_n94) );
  INV_X1 my_filter_adder_mult_7_multiplication_mult_21_U211 ( .A(
        my_filter_q_reg_chain_8__4_), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_n95) );
  INV_X1 my_filter_adder_mult_7_multiplication_mult_21_U210 ( .A(
        my_filter_q_reg_chain_8__2_), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_n97) );
  INV_X1 my_filter_adder_mult_7_multiplication_mult_21_U209 ( .A(
        my_filter_q_reg_chain_8__3_), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_n96) );
  AND2_X1 my_filter_adder_mult_7_multiplication_mult_21_U208 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_13__12_), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_13__13_), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_n3) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U207 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n100), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_13__13_) );
  AND2_X1 my_filter_adder_mult_7_multiplication_mult_21_U206 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_13__9_), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_13__10_), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_n51) );
  AND2_X1 my_filter_adder_mult_7_multiplication_mult_21_U205 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_13__7_), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_13__8_), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_n50) );
  AND2_X1 my_filter_adder_mult_7_multiplication_mult_21_U204 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_13__10_), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_13__11_), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_n48) );
  AND2_X1 my_filter_adder_mult_7_multiplication_mult_21_U203 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_13__8_), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_13__9_), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_n47) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U202 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_12__11_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U201 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_12__10_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U200 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_11__11_) );
  AND2_X1 my_filter_adder_mult_7_multiplication_mult_21_U199 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_13__5_), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_13__6_), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_n44) );
  AND2_X1 my_filter_adder_mult_7_multiplication_mult_21_U198 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_13__3_), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_13__4_), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_n36) );
  AND2_X1 my_filter_adder_mult_7_multiplication_mult_21_U197 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_13__1_), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_13__2_), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_n43) );
  AND2_X1 my_filter_adder_mult_7_multiplication_mult_21_U196 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_13__6_), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_13__7_), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_n42) );
  AND2_X1 my_filter_adder_mult_7_multiplication_mult_21_U195 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_13__4_), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_13__5_), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_n41) );
  AND2_X1 my_filter_adder_mult_7_multiplication_mult_21_U194 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_13__2_), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_13__3_), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_n40) );
  AND2_X1 my_filter_adder_mult_7_multiplication_mult_21_U193 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_13__0_), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_13__1_), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_n35) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U192 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_12__1_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U191 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_10__0_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U190 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_11__0_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U189 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_11__1_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U188 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_10__1_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U187 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_8__0_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U186 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n113), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_9__0_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U185 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n112), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_9__1_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U184 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n110), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_9__3_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U183 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_8__1_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U182 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_8__3_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U181 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_6__0_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U180 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_7__0_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U179 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_7__1_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U178 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_7__3_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U177 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_7__4_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U176 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_7__5_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U175 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_6__1_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U174 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_6__3_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U173 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_6__5_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U172 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_4__0_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U171 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_5__0_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U170 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_5__1_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U169 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_5__3_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U168 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_5__4_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U167 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_5__5_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U166 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_5__6_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U165 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_4__1_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U164 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_4__3_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U163 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_4__5_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U162 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_2__0_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U161 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_3__0_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U160 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_3__1_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U159 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_3__3_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U158 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_3__4_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U157 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_3__5_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U156 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_3__6_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U155 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_3__7_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U154 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_12__9_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U153 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_11__10_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U152 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_12__7_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U151 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_12__8_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U150 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_10__11_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U149 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_11__8_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U148 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_11__9_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U147 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_12__5_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U146 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_12__6_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U145 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_10__9_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U144 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_10__10_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U143 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_11__6_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U142 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_11__7_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U141 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n103), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_9__10_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U140 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n102), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_9__11_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U139 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_12__2_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U138 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_12__3_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U137 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_12__4_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U136 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_10__7_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U135 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_10__8_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U134 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_8__11_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U133 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_11__3_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U132 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_11__4_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U131 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_11__5_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U130 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n105), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_9__8_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U129 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n104), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_9__9_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U128 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_10__4_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U127 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_10__5_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U126 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_10__6_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U125 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_8__9_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U124 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_8__10_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U123 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_11__2_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U122 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n108), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_9__5_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U121 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n107), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_9__6_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U120 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n106), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_9__7_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U119 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_7__10_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U118 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_7__11_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U117 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_10__2_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U116 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_10__3_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U115 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_8__6_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U114 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_8__7_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U113 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_8__8_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U112 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_6__11_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U111 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n111), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_9__2_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U110 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n109), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_9__4_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U109 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_7__7_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U108 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_7__8_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U107 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_7__9_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U106 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_8__2_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U105 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_8__4_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U104 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_8__5_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U103 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_6__8_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U102 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_6__9_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U101 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_6__10_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U100 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_7__2_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U99 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_7__6_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U98 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_5__9_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U97 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_5__10_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U96 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_5__11_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U95 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_6__2_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U94 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_6__4_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U93 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_6__6_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U92 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_6__7_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U91 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_4__10_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U90 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_4__11_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U89 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_5__2_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U88 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_5__7_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U87 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_5__8_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U86 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_3__11_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U85 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_4__2_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U84 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_4__4_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U83 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_4__6_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U82 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_4__7_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U81 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_4__8_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U80 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_4__9_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U79 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_3__2_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U78 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_3__8_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U77 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_3__9_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U76 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_3__10_) );
  AND2_X1 my_filter_adder_mult_7_multiplication_mult_21_U75 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_ab_0__2_), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_ab_1__1_), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_n14) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U74 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_2__1_) );
  AND2_X1 my_filter_adder_mult_7_multiplication_mult_21_U73 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_ab_0__3_), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_ab_1__2_), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_n13) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U72 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_2__2_) );
  AND2_X1 my_filter_adder_mult_7_multiplication_mult_21_U71 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_ab_0__4_), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_ab_1__3_), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_n12) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U70 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_2__3_) );
  AND2_X1 my_filter_adder_mult_7_multiplication_mult_21_U69 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_ab_0__5_), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_ab_1__4_), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_n11) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U68 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_2__4_) );
  AND2_X1 my_filter_adder_mult_7_multiplication_mult_21_U67 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_ab_0__6_), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_ab_1__5_), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_n10) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U66 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_2__5_) );
  AND2_X1 my_filter_adder_mult_7_multiplication_mult_21_U65 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_ab_0__7_), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_ab_1__6_), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_n9) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U64 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_2__6_) );
  AND2_X1 my_filter_adder_mult_7_multiplication_mult_21_U63 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_ab_0__8_), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_ab_1__7_), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_n8) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U62 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_2__7_) );
  AND2_X1 my_filter_adder_mult_7_multiplication_mult_21_U61 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_ab_0__9_), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_ab_1__8_), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_n7) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U60 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_2__8_) );
  AND2_X1 my_filter_adder_mult_7_multiplication_mult_21_U59 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_ab_0__10_), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_ab_1__9_), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_n6) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U58 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_2__9_) );
  AND2_X1 my_filter_adder_mult_7_multiplication_mult_21_U57 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_ab_0__11_), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_ab_1__10_), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_n5) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U56 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_2__10_) );
  AND2_X1 my_filter_adder_mult_7_multiplication_mult_21_U55 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_ab_0__12_), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_ab_1__11_), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_n4) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U54 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_2__11_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U52 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_1__12_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U51 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_1__2_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U50 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_1__3_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U48 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_1__4_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U47 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_1__5_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U44 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_1__6_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U43 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_1__7_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U42 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_1__8_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U41 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_1__9_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U40 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_1__10_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U36 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_1__11_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U35 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_0__2_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U14 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_0__3_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U13 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_0__4_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U12 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_0__5_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U11 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_0__6_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U10 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_0__7_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U9 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_0__8_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U8 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_0__9_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U7 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_0__10_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U6 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_0__11_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U5 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_0__12_) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U4 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n98), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n112), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_ab_1__1_) );
  AND2_X1 my_filter_adder_mult_7_multiplication_mult_21_U3 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_13__11_), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_13__12_), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_n52) );
  INV_X1 my_filter_adder_mult_7_multiplication_mult_21_U2 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_13__13_), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_n85) );
  XOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U49 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_13__10_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_13__11_), .Z(
        my_filter_adder_mult_7_multiplication_mult_21_n49) );
  XOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U46 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_13__11_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_13__12_), .Z(
        my_filter_adder_mult_7_multiplication_mult_21_n46) );
  XOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U45 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_13__9_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_13__10_), .Z(
        my_filter_adder_mult_7_multiplication_mult_21_n45) );
  XOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U39 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_13__5_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_13__6_), .Z(
        my_filter_adder_mult_7_multiplication_mult_21_n39) );
  XOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U38 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_13__3_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_13__4_), .Z(
        my_filter_adder_mult_7_multiplication_mult_21_n38) );
  XOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U37 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_13__1_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_13__2_), .Z(
        my_filter_adder_mult_7_multiplication_mult_21_n37) );
  XOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U34 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_13__8_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_13__9_), .Z(
        my_filter_adder_mult_7_multiplication_mult_21_n34) );
  XOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U33 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_13__6_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_13__7_), .Z(
        my_filter_adder_mult_7_multiplication_mult_21_n33) );
  XOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U32 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_13__7_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_13__8_), .Z(
        my_filter_adder_mult_7_multiplication_mult_21_n32) );
  XOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U31 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_13__4_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_13__5_), .Z(
        my_filter_adder_mult_7_multiplication_mult_21_n31) );
  XOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U30 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_13__2_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_13__3_), .Z(
        my_filter_adder_mult_7_multiplication_mult_21_n30) );
  XOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U29 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_13__0_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_13__1_), .Z(
        my_filter_adder_mult_7_multiplication_mult_21_n29) );
  XOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U27 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_1__1_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_ab_0__2_), .Z(
        my_filter_adder_mult_7_multiplication_mult_21_n28) );
  XOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U26 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_13__12_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_13__13_), .Z(
        my_filter_adder_mult_7_multiplication_mult_21_n27) );
  XOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U25 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_1__12_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_ab_0__13_), .Z(
        my_filter_adder_mult_7_multiplication_mult_21_n26) );
  XOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U24 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_1__2_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_ab_0__3_), .Z(
        my_filter_adder_mult_7_multiplication_mult_21_n25) );
  XOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U23 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_1__3_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_ab_0__4_), .Z(
        my_filter_adder_mult_7_multiplication_mult_21_n24) );
  XOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U22 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_1__4_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_ab_0__5_), .Z(
        my_filter_adder_mult_7_multiplication_mult_21_n23) );
  XOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U21 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_1__5_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_ab_0__6_), .Z(
        my_filter_adder_mult_7_multiplication_mult_21_n22) );
  XOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U20 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_1__6_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_ab_0__7_), .Z(
        my_filter_adder_mult_7_multiplication_mult_21_n21) );
  XOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U19 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_1__7_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_ab_0__8_), .Z(
        my_filter_adder_mult_7_multiplication_mult_21_n20) );
  XOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U18 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_1__8_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_ab_0__9_), .Z(
        my_filter_adder_mult_7_multiplication_mult_21_n19) );
  XOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U17 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_1__9_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_ab_0__10_), .Z(
        my_filter_adder_mult_7_multiplication_mult_21_n18) );
  XOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U16 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_1__10_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_ab_0__11_), .Z(
        my_filter_adder_mult_7_multiplication_mult_21_n17) );
  XOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_U15 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_1__11_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_ab_0__12_), .Z(
        my_filter_adder_mult_7_multiplication_mult_21_n16) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S3_2_12 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_2__12_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_n15), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_ab_1__13_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_2__12_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_2__12_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_2_11 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_2__11_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_n4), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_n26), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_2__11_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_2__11_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_2_10 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_2__10_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_n5), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_n16), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_2__10_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_2__10_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_2_9 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_2__9_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_n6), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_n17), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_2__9_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_2__9_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_2_8 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_2__8_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_n7), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_n18), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_2__8_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_2__8_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_2_7 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_2__7_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_n8), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_n19), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_2__7_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_2__7_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_2_6 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_2__6_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_n9), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_n20), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_2__6_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_2__6_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_2_5 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_2__5_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_n10), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_n21), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_2__5_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_2__5_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_2_4 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_2__4_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_n11), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_n22), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_2__4_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_2__4_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_2_3 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_2__3_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_n12), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_n23), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_2__3_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_2__3_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_2_2 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_2__2_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_n13), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_n24), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_2__2_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_2__2_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_2_1 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_2__1_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_n14), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_n25), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_2__1_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_2__1_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S1_2_0 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_2__0_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_1__0_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_n28), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_2__0_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_A1_0_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S3_3_12 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_3__12_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_2__12_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_ab_2__13_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_3__12_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_3__12_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_3_11 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_3__11_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_2__11_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_2__12_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_3__11_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_3__11_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_3_10 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_3__10_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_2__10_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_2__11_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_3__10_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_3__10_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_3_9 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_3__9_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_2__9_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_2__10_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_3__9_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_3__9_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_3_8 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_3__8_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_2__8_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_2__9_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_3__8_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_3__8_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_3_7 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_3__7_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_2__7_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_2__8_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_3__7_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_3__7_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_3_6 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_3__6_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_2__6_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_2__7_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_3__6_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_3__6_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_3_5 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_3__5_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_2__5_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_2__6_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_3__5_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_3__5_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_3_4 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_3__4_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_2__4_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_2__5_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_3__4_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_3__4_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_3_3 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_3__3_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_2__3_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_2__4_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_3__3_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_3__3_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_3_2 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_3__2_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_2__2_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_2__3_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_3__2_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_3__2_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_3_1 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_3__1_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_2__1_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_2__2_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_3__1_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_3__1_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S1_3_0 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_3__0_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_2__0_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_2__1_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_3__0_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_A1_1_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S3_4_12 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_4__12_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_3__12_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_ab_3__13_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_4__12_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_4__12_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_4_11 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_4__11_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_3__11_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_3__12_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_4__11_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_4__11_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_4_10 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_4__10_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_3__10_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_3__11_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_4__10_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_4__10_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_4_9 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_4__9_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_3__9_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_3__10_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_4__9_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_4__9_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_4_8 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_4__8_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_3__8_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_3__9_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_4__8_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_4__8_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_4_7 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_4__7_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_3__7_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_3__8_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_4__7_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_4__7_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_4_6 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_4__6_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_3__6_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_3__7_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_4__6_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_4__6_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_4_5 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_4__5_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_3__5_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_3__6_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_4__5_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_4__5_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_4_4 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_4__4_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_3__4_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_3__5_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_4__4_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_4__4_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_4_3 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_4__3_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_3__3_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_3__4_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_4__3_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_4__3_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_4_2 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_4__2_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_3__2_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_3__3_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_4__2_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_4__2_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_4_1 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_4__1_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_3__1_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_3__2_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_4__1_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_4__1_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S1_4_0 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_4__0_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_3__0_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_3__1_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_4__0_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_A1_2_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S3_5_12 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_5__12_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_4__12_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_ab_4__13_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_5__12_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_5__12_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_5_11 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_5__11_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_4__11_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_4__12_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_5__11_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_5__11_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_5_10 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_5__10_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_4__10_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_4__11_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_5__10_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_5__10_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_5_9 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_5__9_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_4__9_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_4__10_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_5__9_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_5__9_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_5_8 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_5__8_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_4__8_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_4__9_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_5__8_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_5__8_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_5_7 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_5__7_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_4__7_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_4__8_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_5__7_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_5__7_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_5_6 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_5__6_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_4__6_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_4__7_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_5__6_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_5__6_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_5_5 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_5__5_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_4__5_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_4__6_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_5__5_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_5__5_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_5_4 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_5__4_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_4__4_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_4__5_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_5__4_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_5__4_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_5_3 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_5__3_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_4__3_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_4__4_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_5__3_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_5__3_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_5_2 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_5__2_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_4__2_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_4__3_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_5__2_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_5__2_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_5_1 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_5__1_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_4__1_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_4__2_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_5__1_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_5__1_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S1_5_0 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_5__0_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_4__0_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_4__1_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_5__0_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_A1_3_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S3_6_12 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_6__12_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_5__12_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_ab_5__13_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_6__12_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_6__12_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_6_11 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_6__11_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_5__11_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_5__12_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_6__11_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_6__11_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_6_10 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_6__10_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_5__10_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_5__11_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_6__10_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_6__10_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_6_9 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_6__9_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_5__9_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_5__10_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_6__9_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_6__9_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_6_8 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_6__8_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_5__8_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_5__9_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_6__8_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_6__8_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_6_7 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_6__7_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_5__7_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_5__8_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_6__7_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_6__7_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_6_6 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_6__6_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_5__6_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_5__7_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_6__6_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_6__6_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_6_5 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_6__5_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_5__5_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_5__6_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_6__5_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_6__5_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_6_4 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_6__4_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_5__4_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_5__5_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_6__4_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_6__4_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_6_3 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_6__3_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_5__3_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_5__4_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_6__3_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_6__3_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_6_2 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_6__2_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_5__2_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_5__3_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_6__2_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_6__2_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_6_1 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_6__1_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_5__1_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_5__2_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_6__1_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_6__1_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S1_6_0 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_6__0_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_5__0_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_5__1_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_6__0_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_A1_4_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S3_7_12 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_7__12_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_6__12_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_ab_6__13_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_7__12_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_7__12_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_7_11 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_7__11_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_6__11_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_6__12_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_7__11_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_7__11_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_7_10 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_7__10_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_6__10_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_6__11_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_7__10_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_7__10_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_7_9 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_7__9_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_6__9_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_6__10_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_7__9_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_7__9_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_7_8 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_7__8_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_6__8_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_6__9_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_7__8_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_7__8_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_7_7 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_7__7_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_6__7_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_6__8_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_7__7_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_7__7_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_7_6 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_7__6_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_6__6_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_6__7_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_7__6_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_7__6_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_7_5 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_7__5_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_6__5_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_6__6_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_7__5_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_7__5_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_7_4 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_7__4_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_6__4_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_6__5_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_7__4_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_7__4_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_7_3 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_7__3_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_6__3_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_6__4_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_7__3_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_7__3_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_7_2 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_7__2_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_6__2_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_6__3_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_7__2_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_7__2_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_7_1 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_7__1_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_6__1_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_6__2_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_7__1_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_7__1_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S1_7_0 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_7__0_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_6__0_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_6__1_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_7__0_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_A1_5_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S3_8_12 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_8__12_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_7__12_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_ab_7__13_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_8__12_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_8__12_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_8_11 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_8__11_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_7__11_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_7__12_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_8__11_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_8__11_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_8_10 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_8__10_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_7__10_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_7__11_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_8__10_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_8__10_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_8_9 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_8__9_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_7__9_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_7__10_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_8__9_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_8__9_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_8_8 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_8__8_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_7__8_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_7__9_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_8__8_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_8__8_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_8_7 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_8__7_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_7__7_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_7__8_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_8__7_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_8__7_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_8_6 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_8__6_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_7__6_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_7__7_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_8__6_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_8__6_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_8_5 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_8__5_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_7__5_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_7__6_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_8__5_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_8__5_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_8_4 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_8__4_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_7__4_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_7__5_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_8__4_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_8__4_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_8_3 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_8__3_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_7__3_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_7__4_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_8__3_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_8__3_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_8_2 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_8__2_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_7__2_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_7__3_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_8__2_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_8__2_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_8_1 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_8__1_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_7__1_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_7__2_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_8__1_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_8__1_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S1_8_0 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_8__0_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_7__0_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_7__1_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_8__0_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_A1_6_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S3_9_12 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_9__12_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_8__12_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_ab_8__13_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_9__12_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_9__12_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_9_11 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_9__11_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_8__11_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_8__12_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_9__11_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_9__11_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_9_10 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_9__10_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_8__10_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_8__11_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_9__10_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_9__10_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_9_9 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_9__9_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_8__9_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_8__10_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_9__9_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_9__9_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_9_8 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_9__8_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_8__8_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_8__9_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_9__8_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_9__8_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_9_7 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_9__7_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_8__7_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_8__8_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_9__7_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_9__7_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_9_6 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_9__6_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_8__6_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_8__7_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_9__6_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_9__6_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_9_5 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_9__5_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_8__5_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_8__6_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_9__5_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_9__5_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_9_4 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_9__4_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_8__4_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_8__5_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_9__4_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_9__4_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_9_3 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_9__3_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_8__3_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_8__4_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_9__3_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_9__3_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_9_2 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_9__2_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_8__2_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_8__3_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_9__2_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_9__2_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_9_1 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_9__1_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_8__1_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_8__2_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_9__1_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_9__1_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S1_9_0 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_9__0_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_8__0_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_8__1_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_9__0_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_A1_7_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S3_10_12 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_10__12_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_9__12_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_ab_9__13_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_10__12_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_10__12_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_10_11 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_10__11_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_9__11_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_9__12_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_10__11_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_10__11_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_10_10 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_10__10_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_9__10_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_9__11_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_10__10_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_10__10_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_10_9 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_10__9_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_9__9_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_9__10_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_10__9_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_10__9_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_10_8 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_10__8_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_9__8_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_9__9_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_10__8_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_10__8_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_10_7 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_10__7_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_9__7_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_9__8_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_10__7_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_10__7_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_10_6 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_10__6_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_9__6_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_9__7_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_10__6_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_10__6_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_10_5 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_10__5_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_9__5_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_9__6_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_10__5_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_10__5_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_10_4 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_10__4_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_9__4_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_9__5_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_10__4_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_10__4_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_10_3 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_10__3_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_9__3_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_9__4_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_10__3_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_10__3_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_10_2 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_10__2_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_9__2_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_9__3_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_10__2_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_10__2_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_10_1 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_10__1_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_9__1_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_9__2_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_10__1_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_10__1_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S1_10_0 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_10__0_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_9__0_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_9__1_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_10__0_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_A1_8_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S3_11_12 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_11__12_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_10__12_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_ab_10__13_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_11__12_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_11__12_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_11_11 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_11__11_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_10__11_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_10__12_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_11__11_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_11__11_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_11_10 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_11__10_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_10__10_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_10__11_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_11__10_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_11__10_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_11_9 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_11__9_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_10__9_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_10__10_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_11__9_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_11__9_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_11_8 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_11__8_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_10__8_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_10__9_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_11__8_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_11__8_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_11_7 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_11__7_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_10__7_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_10__8_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_11__7_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_11__7_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_11_6 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_11__6_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_10__6_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_10__7_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_11__6_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_11__6_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_11_5 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_11__5_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_10__5_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_10__6_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_11__5_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_11__5_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_11_4 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_11__4_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_10__4_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_10__5_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_11__4_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_11__4_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_11_3 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_11__3_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_10__3_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_10__4_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_11__3_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_11__3_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_11_2 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_11__2_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_10__2_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_10__3_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_11__2_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_11__2_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_11_1 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_11__1_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_10__1_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_10__2_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_11__1_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_11__1_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S1_11_0 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_11__0_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_10__0_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_10__1_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_11__0_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_A1_9_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S3_12_12 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_12__12_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_11__12_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_ab_11__13_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_12__12_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_12__12_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_12_11 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_12__11_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_11__11_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_11__12_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_12__11_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_12__11_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_12_10 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_12__10_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_11__10_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_11__11_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_12__10_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_12__10_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_12_9 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_12__9_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_11__9_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_11__10_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_12__9_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_12__9_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_12_8 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_12__8_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_11__8_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_11__9_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_12__8_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_12__8_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_12_7 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_12__7_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_11__7_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_11__8_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_12__7_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_12__7_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_12_6 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_12__6_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_11__6_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_11__7_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_12__6_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_12__6_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_12_5 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_12__5_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_11__5_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_11__6_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_12__5_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_12__5_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_12_4 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_12__4_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_11__4_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_11__5_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_12__4_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_12__4_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_12_3 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_12__3_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_11__3_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_11__4_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_12__3_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_12__3_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_12_2 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_12__2_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_11__2_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_11__3_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_12__2_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_12__2_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S2_12_1 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_12__1_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_11__1_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_11__2_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_12__1_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_12__1_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S1_12_0 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_12__0_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_11__0_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_11__1_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_12__0_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_A1_10_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S14_13 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_n86), .B(
        my_filter_adder_mult_7_multiplication_mult_21_n100), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_ab_13__13_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_13__13_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_13__13_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S5_12 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_13__12_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_12__12_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_ab_12__13_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_13__12_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_13__12_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S4_11 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_13__11_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_12__11_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_12__12_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_13__11_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_13__11_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S4_10 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_13__10_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_12__10_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_12__11_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_13__10_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_13__10_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S4_9 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_13__9_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_12__9_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_12__10_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_13__9_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_13__9_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S4_8 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_13__8_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_12__8_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_12__9_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_13__8_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_13__8_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S4_7 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_13__7_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_12__7_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_12__8_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_13__7_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_13__7_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S4_6 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_13__6_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_12__6_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_12__7_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_13__6_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_13__6_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S4_5 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_13__5_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_12__5_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_12__6_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_13__5_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_13__5_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S4_4 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_13__4_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_12__4_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_12__5_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_13__4_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_13__4_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S4_3 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_13__3_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_12__3_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_12__4_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_13__3_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_13__3_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S4_2 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_13__2_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_12__2_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_12__3_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_13__2_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_13__2_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S4_1 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_13__1_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_12__1_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_12__2_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_13__1_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_13__1_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S4_0 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_ab_13__0_), .B(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_12__0_), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_12__1_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_CARRYB_13__0_), .S(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_13__0_) );
  FA_X1 my_filter_adder_mult_7_multiplication_mult_21_S14_13_0 ( .A(
        my_filter_q_reg_chain_8__13_), .B(my_filter_q_reg_coeff[41]), .CI(
        my_filter_adder_mult_7_multiplication_mult_21_SUMB_13__0_), .CO(
        my_filter_adder_mult_7_multiplication_mult_21_A2_12_), .S(
        my_filter_adder_mult_7_res_mult[0]) );
  NAND2_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U72 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_A2_12_), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n29), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n56) );
  OAI21_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U71 ( .B1(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n15), .B2(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n16), .A(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n17), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n13) );
  OAI21_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U70 ( .B1(
        my_filter_adder_mult_7_multiplication_mult_21_A2_12_), .B2(
        my_filter_adder_mult_7_multiplication_mult_21_n29), .A(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n56), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n59) );
  INV_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U69 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n59), .ZN(
        my_filter_adder_mult_7_res_mult[1]) );
  AND2_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U68 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n51), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n49), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n20) );
  AND2_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U66 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n50), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n34), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n28) );
  NAND2_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U65 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n48), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n46), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n17) );
  NAND2_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U64 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n47), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n45), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n25) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U63 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n48), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n46), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n15) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U61 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n47), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n45), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n23) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U60 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n51), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n49), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n21) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U59 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n50), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n34), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n29) );
  AND2_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U58 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n44), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n33), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n36) );
  AND2_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U56 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n36), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n31), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n44) );
  AND2_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U55 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n43), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n30), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n52) );
  NAND2_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U54 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n42), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n32), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n33) );
  NAND2_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U53 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n41), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n39), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n41) );
  NAND2_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U51 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n40), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n38), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n49) );
  NAND2_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U50 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n35), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n37), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n57) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U49 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n42), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n32), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n31) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U48 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n41), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n39), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n39) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U46 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n40), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n38), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n47) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U45 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n35), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n37), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n55) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U44 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n44), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n33), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n37) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U43 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n36), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n31), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n45) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U41 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_n43), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_n30), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n53) );
  OAI21_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U40 ( .B1(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n55), .B2(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n56), .A(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n57), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n51) );
  INV_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U39 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n55), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n60) );
  NAND2_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U38 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n60), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n57), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n58) );
  OAI21_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U36 ( .B1(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n23), .B2(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n24), .A(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n25), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n19) );
  OAI21_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U35 ( .B1(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n31), .B2(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n32), .A(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n33), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n27) );
  OAI21_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U34 ( .B1(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n39), .B2(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n40), .A(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n41), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n35) );
  OAI21_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U33 ( .B1(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n47), .B2(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n48), .A(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n49), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n43) );
  INV_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U31 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n21), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n63) );
  AOI21_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U30 ( .B1(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n63), .B2(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n19), .A(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n20), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n16) );
  INV_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U29 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n29), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n71) );
  AOI21_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U28 ( .B1(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n71), .B2(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n27), .A(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n28), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n24) );
  INV_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U26 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n37), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n69) );
  AOI21_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U25 ( .B1(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n69), .B2(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n35), .A(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n36), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n32) );
  INV_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U24 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n45), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n67) );
  AOI21_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U23 ( .B1(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n67), .B2(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n43), .A(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n44), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n40) );
  INV_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U21 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n53), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n65) );
  AOI21_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U20 ( .B1(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n65), .B2(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n51), .A(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n52), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n48) );
  INV_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U19 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n15), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n62) );
  NAND2_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U18 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n62), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n17), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n18) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U16 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n20), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n21), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n22) );
  INV_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U13 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n23), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n64) );
  NAND2_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U12 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n64), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n25), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n26) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U11 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n28), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n29), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n30) );
  INV_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U10 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n31), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n70) );
  NAND2_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U9 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n70), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n33), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n34) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U8 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n36), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n37), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n38) );
  INV_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U7 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n39), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n68) );
  NAND2_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U6 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n68), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n41), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n42) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U5 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n44), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n45), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n46) );
  INV_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U4 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n47), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n66) );
  NAND2_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U3 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n66), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n49), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n50) );
  NOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U2 ( .A1(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n52), .A2(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n53), .ZN(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n54) );
  XOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U67 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n56), .B(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n58), .Z(
        my_filter_adder_mult_7_res_mult[2]) );
  XOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U62 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n51), .B(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n54), .Z(
        my_filter_adder_mult_7_res_mult[3]) );
  XOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U57 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n50), .B(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n48), .Z(
        my_filter_adder_mult_7_res_mult[4]) );
  XOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U52 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n43), .B(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n46), .Z(
        my_filter_adder_mult_7_res_mult[5]) );
  XOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U47 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n42), .B(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n40), .Z(
        my_filter_adder_mult_7_res_mult[6]) );
  XOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U42 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n35), .B(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n38), .Z(
        my_filter_adder_mult_7_res_mult[7]) );
  XOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U37 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n34), .B(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n32), .Z(
        my_filter_adder_mult_7_res_mult[8]) );
  XOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U32 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n27), .B(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n30), .Z(
        my_filter_adder_mult_7_res_mult[9]) );
  XOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U27 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n26), .B(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n24), .Z(
        my_filter_adder_mult_7_res_mult[10]) );
  XOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U22 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n19), .B(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n22), .Z(
        my_filter_adder_mult_7_res_mult[11]) );
  XOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U17 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n18), .B(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n16), .Z(
        my_filter_adder_mult_7_res_mult[12]) );
  XOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U15 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_n52), .B(
        my_filter_adder_mult_7_multiplication_mult_21_n27), .Z(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n14) );
  XOR2_X1 my_filter_adder_mult_7_multiplication_mult_21_FS_1_U14 ( .A(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n13), .B(
        my_filter_adder_mult_7_multiplication_mult_21_FS_1_n14), .Z(
        my_filter_adder_mult_7_res_mult[13]) );
  AND2_X1 my_filter_adder_mult_7_addition_add_19_U1 ( .A1(
        my_filter_data_sum[42]), .A2(my_filter_adder_mult_7_res_mult[0]), .ZN(
        my_filter_adder_mult_7_addition_add_19_n1) );
  XOR2_X1 my_filter_adder_mult_7_addition_add_19_U2 ( .A(
        my_filter_data_sum[42]), .B(my_filter_adder_mult_7_res_mult[0]), .Z(
        my_filter_data_sum[28]) );
  FA_X1 my_filter_adder_mult_7_addition_add_19_U1_1 ( .A(
        my_filter_adder_mult_7_res_mult[1]), .B(my_filter_data_sum[43]), .CI(
        my_filter_adder_mult_7_addition_add_19_n1), .CO(
        my_filter_adder_mult_7_addition_add_19_carry[2]), .S(
        my_filter_data_sum[29]) );
  FA_X1 my_filter_adder_mult_7_addition_add_19_U1_2 ( .A(
        my_filter_adder_mult_7_res_mult[2]), .B(my_filter_data_sum[44]), .CI(
        my_filter_adder_mult_7_addition_add_19_carry[2]), .CO(
        my_filter_adder_mult_7_addition_add_19_carry[3]), .S(
        my_filter_data_sum[30]) );
  FA_X1 my_filter_adder_mult_7_addition_add_19_U1_3 ( .A(
        my_filter_adder_mult_7_res_mult[3]), .B(my_filter_data_sum[45]), .CI(
        my_filter_adder_mult_7_addition_add_19_carry[3]), .CO(
        my_filter_adder_mult_7_addition_add_19_carry[4]), .S(
        my_filter_data_sum[31]) );
  FA_X1 my_filter_adder_mult_7_addition_add_19_U1_4 ( .A(
        my_filter_adder_mult_7_res_mult[4]), .B(my_filter_data_sum[46]), .CI(
        my_filter_adder_mult_7_addition_add_19_carry[4]), .CO(
        my_filter_adder_mult_7_addition_add_19_carry[5]), .S(
        my_filter_data_sum[32]) );
  FA_X1 my_filter_adder_mult_7_addition_add_19_U1_5 ( .A(
        my_filter_adder_mult_7_res_mult[5]), .B(my_filter_data_sum[47]), .CI(
        my_filter_adder_mult_7_addition_add_19_carry[5]), .CO(
        my_filter_adder_mult_7_addition_add_19_carry[6]), .S(
        my_filter_data_sum[33]) );
  FA_X1 my_filter_adder_mult_7_addition_add_19_U1_6 ( .A(
        my_filter_adder_mult_7_res_mult[6]), .B(my_filter_data_sum[48]), .CI(
        my_filter_adder_mult_7_addition_add_19_carry[6]), .CO(
        my_filter_adder_mult_7_addition_add_19_carry[7]), .S(
        my_filter_data_sum[34]) );
  FA_X1 my_filter_adder_mult_7_addition_add_19_U1_7 ( .A(
        my_filter_adder_mult_7_res_mult[7]), .B(my_filter_data_sum[49]), .CI(
        my_filter_adder_mult_7_addition_add_19_carry[7]), .CO(
        my_filter_adder_mult_7_addition_add_19_carry[8]), .S(
        my_filter_data_sum[35]) );
  FA_X1 my_filter_adder_mult_7_addition_add_19_U1_8 ( .A(
        my_filter_adder_mult_7_res_mult[8]), .B(my_filter_data_sum[50]), .CI(
        my_filter_adder_mult_7_addition_add_19_carry[8]), .CO(
        my_filter_adder_mult_7_addition_add_19_carry[9]), .S(
        my_filter_data_sum[36]) );
  FA_X1 my_filter_adder_mult_7_addition_add_19_U1_9 ( .A(
        my_filter_adder_mult_7_res_mult[9]), .B(my_filter_data_sum[51]), .CI(
        my_filter_adder_mult_7_addition_add_19_carry[9]), .CO(
        my_filter_adder_mult_7_addition_add_19_carry[10]), .S(
        my_filter_data_sum[37]) );
  FA_X1 my_filter_adder_mult_7_addition_add_19_U1_10 ( .A(
        my_filter_adder_mult_7_res_mult[10]), .B(my_filter_data_sum[52]), .CI(
        my_filter_adder_mult_7_addition_add_19_carry[10]), .CO(
        my_filter_adder_mult_7_addition_add_19_carry[11]), .S(
        my_filter_data_sum[38]) );
  FA_X1 my_filter_adder_mult_7_addition_add_19_U1_11 ( .A(
        my_filter_adder_mult_7_res_mult[11]), .B(my_filter_data_sum[53]), .CI(
        my_filter_adder_mult_7_addition_add_19_carry[11]), .CO(
        my_filter_adder_mult_7_addition_add_19_carry[12]), .S(
        my_filter_data_sum[39]) );
  FA_X1 my_filter_adder_mult_7_addition_add_19_U1_12 ( .A(
        my_filter_adder_mult_7_res_mult[12]), .B(my_filter_data_sum[54]), .CI(
        my_filter_adder_mult_7_addition_add_19_carry[12]), .CO(
        my_filter_adder_mult_7_addition_add_19_carry[13]), .S(
        my_filter_data_sum[40]) );
  FA_X1 my_filter_adder_mult_7_addition_add_19_U1_13 ( .A(
        my_filter_adder_mult_7_res_mult[13]), .B(my_filter_data_sum[55]), .CI(
        my_filter_adder_mult_7_addition_add_19_carry[13]), .S(
        my_filter_data_sum[41]) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U276 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_12__12_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U275 ( .A1(
        my_filter_q_reg_chain_9__11_), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_11__13_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U274 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_11__12_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U273 ( .A1(
        my_filter_q_reg_chain_9__10_), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_10__13_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U272 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_10__12_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U271 ( .A1(
        my_filter_q_reg_chain_9__9_), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_9__13_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U270 ( .A1(
        my_filter_q_reg_chain_9__8_), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_8__13_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U269 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n101), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_9__12_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U268 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_8__12_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U267 ( .A1(
        my_filter_q_reg_chain_9__7_), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_7__13_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U266 ( .A1(
        my_filter_q_reg_coeff[24]), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_13__10_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U265 ( .A1(
        my_filter_q_reg_coeff[25]), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_13__11_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U264 ( .A1(
        my_filter_q_reg_coeff[22]), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_13__8_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U263 ( .A1(
        my_filter_q_reg_coeff[23]), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_13__9_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U262 ( .A1(
        my_filter_q_reg_coeff[26]), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_13__12_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U261 ( .A1(
        my_filter_q_reg_chain_9__12_), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_12__13_) );
  INV_X1 my_filter_adder_mult_8_multiplication_mult_21_U260 ( .A(
        my_filter_q_reg_chain_9__9_), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_n90) );
  INV_X1 my_filter_adder_mult_8_multiplication_mult_21_U259 ( .A(
        my_filter_q_reg_chain_9__12_), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_n87) );
  INV_X1 my_filter_adder_mult_8_multiplication_mult_21_U258 ( .A(
        my_filter_q_reg_chain_9__11_), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_n88) );
  INV_X1 my_filter_adder_mult_8_multiplication_mult_21_U257 ( .A(
        my_filter_q_reg_chain_9__10_), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_n89) );
  INV_X1 my_filter_adder_mult_8_multiplication_mult_21_U256 ( .A(
        my_filter_q_reg_chain_9__8_), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_n91) );
  INV_X1 my_filter_adder_mult_8_multiplication_mult_21_U255 ( .A(
        my_filter_q_reg_chain_9__7_), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_n92) );
  INV_X1 my_filter_adder_mult_8_multiplication_mult_21_U254 ( .A(
        my_filter_q_reg_chain_9__13_), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_n86) );
  AND2_X1 my_filter_adder_mult_8_multiplication_mult_21_U253 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_ab_0__13_), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_ab_1__12_), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_n15) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U252 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_2__12_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U251 ( .A1(
        my_filter_q_reg_chain_9__1_), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_1__13_) );
  AND3_X1 my_filter_adder_mult_8_multiplication_mult_21_U250 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_ab_1__1_), .A2(
        my_filter_q_reg_coeff[14]), .A3(my_filter_q_reg_chain_9__0_), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_1__0_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U249 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_12__0_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U248 ( .A1(
        my_filter_q_reg_coeff[14]), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_13__0_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U247 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_7__12_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U246 ( .A1(
        my_filter_q_reg_chain_9__6_), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_6__13_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U245 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_6__12_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U244 ( .A1(
        my_filter_q_reg_chain_9__5_), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_5__13_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U243 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_5__12_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U242 ( .A1(
        my_filter_q_reg_chain_9__4_), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_4__13_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U241 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_4__12_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U240 ( .A1(
        my_filter_q_reg_chain_9__3_), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_3__13_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U239 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_3__12_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U238 ( .A1(
        my_filter_q_reg_chain_9__2_), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_2__13_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U237 ( .A1(
        my_filter_q_reg_coeff[20]), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_13__6_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U236 ( .A1(
        my_filter_q_reg_coeff[21]), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_13__7_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U235 ( .A1(
        my_filter_q_reg_coeff[18]), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_13__4_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U234 ( .A1(
        my_filter_q_reg_coeff[19]), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_13__5_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U233 ( .A1(
        my_filter_q_reg_coeff[16]), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_13__2_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U232 ( .A1(
        my_filter_q_reg_coeff[17]), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_13__3_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U231 ( .A1(
        my_filter_q_reg_coeff[15]), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_13__1_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U230 ( .A1(
        my_filter_q_reg_chain_9__0_), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_0__13_) );
  INV_X1 my_filter_adder_mult_8_multiplication_mult_21_U229 ( .A(
        my_filter_q_reg_coeff[27]), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_n100) );
  INV_X1 my_filter_adder_mult_8_multiplication_mult_21_U228 ( .A(
        my_filter_q_reg_coeff[14]), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_n113) );
  INV_X1 my_filter_adder_mult_8_multiplication_mult_21_U227 ( .A(
        my_filter_q_reg_chain_9__0_), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_n99) );
  INV_X1 my_filter_adder_mult_8_multiplication_mult_21_U226 ( .A(
        my_filter_q_reg_coeff[15]), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_n112) );
  INV_X1 my_filter_adder_mult_8_multiplication_mult_21_U225 ( .A(
        my_filter_q_reg_chain_9__1_), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_n98) );
  INV_X1 my_filter_adder_mult_8_multiplication_mult_21_U224 ( .A(
        my_filter_q_reg_coeff[26]), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_n101) );
  INV_X1 my_filter_adder_mult_8_multiplication_mult_21_U223 ( .A(
        my_filter_q_reg_coeff[24]), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_n103) );
  INV_X1 my_filter_adder_mult_8_multiplication_mult_21_U222 ( .A(
        my_filter_q_reg_coeff[25]), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_n102) );
  INV_X1 my_filter_adder_mult_8_multiplication_mult_21_U221 ( .A(
        my_filter_q_reg_coeff[22]), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_n105) );
  INV_X1 my_filter_adder_mult_8_multiplication_mult_21_U220 ( .A(
        my_filter_q_reg_coeff[23]), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_n104) );
  INV_X1 my_filter_adder_mult_8_multiplication_mult_21_U219 ( .A(
        my_filter_q_reg_coeff[20]), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_n107) );
  INV_X1 my_filter_adder_mult_8_multiplication_mult_21_U218 ( .A(
        my_filter_q_reg_coeff[21]), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_n106) );
  INV_X1 my_filter_adder_mult_8_multiplication_mult_21_U217 ( .A(
        my_filter_q_reg_coeff[16]), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_n111) );
  INV_X1 my_filter_adder_mult_8_multiplication_mult_21_U216 ( .A(
        my_filter_q_reg_coeff[17]), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_n110) );
  INV_X1 my_filter_adder_mult_8_multiplication_mult_21_U215 ( .A(
        my_filter_q_reg_coeff[18]), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_n109) );
  INV_X1 my_filter_adder_mult_8_multiplication_mult_21_U214 ( .A(
        my_filter_q_reg_coeff[19]), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_n108) );
  INV_X1 my_filter_adder_mult_8_multiplication_mult_21_U213 ( .A(
        my_filter_q_reg_chain_9__6_), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_n93) );
  INV_X1 my_filter_adder_mult_8_multiplication_mult_21_U212 ( .A(
        my_filter_q_reg_chain_9__5_), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_n94) );
  INV_X1 my_filter_adder_mult_8_multiplication_mult_21_U211 ( .A(
        my_filter_q_reg_chain_9__4_), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_n95) );
  INV_X1 my_filter_adder_mult_8_multiplication_mult_21_U210 ( .A(
        my_filter_q_reg_chain_9__3_), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_n96) );
  INV_X1 my_filter_adder_mult_8_multiplication_mult_21_U209 ( .A(
        my_filter_q_reg_chain_9__2_), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_n97) );
  AND2_X1 my_filter_adder_mult_8_multiplication_mult_21_U208 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_13__12_), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_13__13_), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_n3) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U207 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n100), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_13__13_) );
  AND2_X1 my_filter_adder_mult_8_multiplication_mult_21_U206 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_13__11_), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_13__12_), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_n52) );
  AND2_X1 my_filter_adder_mult_8_multiplication_mult_21_U205 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_13__9_), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_13__10_), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_n50) );
  AND2_X1 my_filter_adder_mult_8_multiplication_mult_21_U204 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_13__7_), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_13__8_), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_n49) );
  AND2_X1 my_filter_adder_mult_8_multiplication_mult_21_U203 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_13__5_), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_13__6_), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_n40) );
  AND2_X1 my_filter_adder_mult_8_multiplication_mult_21_U202 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_13__10_), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_13__11_), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_n47) );
  AND2_X1 my_filter_adder_mult_8_multiplication_mult_21_U201 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_13__8_), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_13__9_), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_n46) );
  AND2_X1 my_filter_adder_mult_8_multiplication_mult_21_U200 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_13__6_), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_13__7_), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_n45) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U199 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_12__11_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U198 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_12__9_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U197 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_12__10_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U196 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_11__10_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U195 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_11__11_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U194 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_10__11_) );
  AND2_X1 my_filter_adder_mult_8_multiplication_mult_21_U193 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_13__3_), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_13__4_), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_n35) );
  AND2_X1 my_filter_adder_mult_8_multiplication_mult_21_U192 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_13__1_), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_13__2_), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_n39) );
  AND2_X1 my_filter_adder_mult_8_multiplication_mult_21_U191 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_13__4_), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_13__5_), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_n34) );
  AND2_X1 my_filter_adder_mult_8_multiplication_mult_21_U190 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_13__2_), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_13__3_), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_n33) );
  AND2_X1 my_filter_adder_mult_8_multiplication_mult_21_U189 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_13__0_), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_13__1_), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_n32) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U188 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_12__1_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U187 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_10__0_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U186 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_11__0_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U185 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_11__1_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U184 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_10__1_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U183 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_8__0_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U182 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n113), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_9__0_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U181 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n112), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_9__1_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U180 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n110), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_9__3_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U179 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_8__1_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U178 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_8__3_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U177 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_6__0_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U176 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_7__0_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U175 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_7__1_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U174 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_7__3_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U173 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_7__4_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U172 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_7__5_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U171 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_6__1_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U170 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_6__3_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U169 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_6__5_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U168 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_4__0_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U167 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_5__0_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U166 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_5__1_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U165 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_5__3_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U164 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_5__4_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U163 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_5__5_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U162 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_5__6_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U161 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_4__1_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U160 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_4__3_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U159 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_4__5_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U158 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_2__0_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U157 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_3__0_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U156 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_3__1_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U155 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_3__3_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U154 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_3__4_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U153 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_3__5_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U152 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_3__6_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U151 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_3__7_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U150 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_12__7_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U149 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_12__8_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U148 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_11__8_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U147 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_11__9_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U146 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_10__9_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U145 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_10__10_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U144 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_12__5_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U143 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_12__6_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U142 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n103), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_9__10_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U141 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n102), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_9__11_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U140 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_11__6_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U139 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_11__7_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U138 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_8__11_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U137 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_10__7_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U136 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_10__8_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U135 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_12__3_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U134 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_12__4_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U133 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n105), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_9__8_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U132 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n104), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_9__9_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U131 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_11__4_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U130 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_11__5_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U129 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_12__2_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U128 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_8__9_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U127 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_8__10_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U126 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_10__5_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U125 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_10__6_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U124 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_11__3_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U123 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_7__10_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U122 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_7__11_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U121 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n107), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_9__6_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U120 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n106), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_9__7_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U119 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_11__2_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U118 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_10__4_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U117 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_6__11_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U116 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_8__7_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U115 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_8__8_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U114 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_10__2_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U113 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_10__3_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U112 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n108), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_9__5_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U111 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_7__8_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U110 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_7__9_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U109 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n111), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_9__2_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U108 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n109), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_9__4_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U107 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_8__6_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U106 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_6__9_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U105 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_6__10_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U104 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_8__2_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U103 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_8__4_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U102 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_8__5_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U101 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_7__7_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U100 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_5__10_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U99 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_5__11_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U98 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_7__2_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U97 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_7__6_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U96 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_6__8_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U95 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_4__11_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U94 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_6__2_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U93 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_6__4_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U92 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_6__6_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U91 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_6__7_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U90 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_5__9_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U89 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_5__2_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U88 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_5__7_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U87 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_5__8_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U86 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_4__10_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U85 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_4__2_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U84 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_4__4_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U83 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_4__6_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U82 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_4__7_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U81 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_4__8_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U80 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_4__9_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U79 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_3__11_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U78 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_3__2_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U77 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_3__8_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U76 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_3__9_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U75 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_3__10_) );
  AND2_X1 my_filter_adder_mult_8_multiplication_mult_21_U74 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_ab_0__2_), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_ab_1__1_), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_n14) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U73 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_2__1_) );
  AND2_X1 my_filter_adder_mult_8_multiplication_mult_21_U72 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_ab_0__3_), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_ab_1__2_), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_n13) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U71 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_2__2_) );
  AND2_X1 my_filter_adder_mult_8_multiplication_mult_21_U70 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_ab_0__4_), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_ab_1__3_), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_n12) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U69 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_2__3_) );
  AND2_X1 my_filter_adder_mult_8_multiplication_mult_21_U68 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_ab_0__5_), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_ab_1__4_), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_n11) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U67 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_2__4_) );
  AND2_X1 my_filter_adder_mult_8_multiplication_mult_21_U66 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_ab_0__6_), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_ab_1__5_), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_n10) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U65 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_2__5_) );
  AND2_X1 my_filter_adder_mult_8_multiplication_mult_21_U64 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_ab_0__7_), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_ab_1__6_), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_n9) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U63 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_2__6_) );
  AND2_X1 my_filter_adder_mult_8_multiplication_mult_21_U62 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_ab_0__8_), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_ab_1__7_), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_n8) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U61 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_2__7_) );
  AND2_X1 my_filter_adder_mult_8_multiplication_mult_21_U60 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_ab_0__9_), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_ab_1__8_), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_n7) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U59 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_2__8_) );
  AND2_X1 my_filter_adder_mult_8_multiplication_mult_21_U58 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_ab_0__10_), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_ab_1__9_), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_n6) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U57 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_2__9_) );
  AND2_X1 my_filter_adder_mult_8_multiplication_mult_21_U56 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_ab_0__11_), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_ab_1__10_), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_n5) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U55 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_2__10_) );
  AND2_X1 my_filter_adder_mult_8_multiplication_mult_21_U54 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_ab_0__12_), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_ab_1__11_), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_n4) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U52 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_2__11_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U50 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_1__12_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U49 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_1__2_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U47 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_1__3_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U46 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_1__4_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U45 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_1__5_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U40 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_1__6_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U39 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_1__7_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U35 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_1__8_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U34 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_1__9_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U33 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_1__10_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U32 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_1__11_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U14 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_0__2_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U13 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_0__3_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U12 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_0__4_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U11 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_0__5_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U10 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_0__6_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U9 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_0__7_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U8 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_0__8_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U7 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_0__9_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U6 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_0__10_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U5 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_0__11_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U4 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_0__12_) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U3 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n98), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n112), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_ab_1__1_) );
  INV_X1 my_filter_adder_mult_8_multiplication_mult_21_U2 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_13__13_), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_n85) );
  XOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U51 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_13__12_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_13__13_), .Z(
        my_filter_adder_mult_8_multiplication_mult_21_n51) );
  XOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U48 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_13__10_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_13__11_), .Z(
        my_filter_adder_mult_8_multiplication_mult_21_n48) );
  XOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U44 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_13__11_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_13__12_), .Z(
        my_filter_adder_mult_8_multiplication_mult_21_n44) );
  XOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U43 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_13__8_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_13__9_), .Z(
        my_filter_adder_mult_8_multiplication_mult_21_n43) );
  XOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U42 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_13__9_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_13__10_), .Z(
        my_filter_adder_mult_8_multiplication_mult_21_n42) );
  XOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U41 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_13__7_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_13__8_), .Z(
        my_filter_adder_mult_8_multiplication_mult_21_n41) );
  XOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U38 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_13__5_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_13__6_), .Z(
        my_filter_adder_mult_8_multiplication_mult_21_n38) );
  XOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U37 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_13__3_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_13__4_), .Z(
        my_filter_adder_mult_8_multiplication_mult_21_n37) );
  XOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U36 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_13__1_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_13__2_), .Z(
        my_filter_adder_mult_8_multiplication_mult_21_n36) );
  XOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U31 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_13__6_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_13__7_), .Z(
        my_filter_adder_mult_8_multiplication_mult_21_n31) );
  XOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U30 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_13__4_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_13__5_), .Z(
        my_filter_adder_mult_8_multiplication_mult_21_n30) );
  XOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U29 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_13__2_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_13__3_), .Z(
        my_filter_adder_mult_8_multiplication_mult_21_n29) );
  XOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U28 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_13__0_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_13__1_), .Z(
        my_filter_adder_mult_8_multiplication_mult_21_n28) );
  XOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U26 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_1__1_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_ab_0__2_), .Z(
        my_filter_adder_mult_8_multiplication_mult_21_n27) );
  XOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U25 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_1__12_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_ab_0__13_), .Z(
        my_filter_adder_mult_8_multiplication_mult_21_n26) );
  XOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U24 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_1__2_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_ab_0__3_), .Z(
        my_filter_adder_mult_8_multiplication_mult_21_n25) );
  XOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U23 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_1__3_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_ab_0__4_), .Z(
        my_filter_adder_mult_8_multiplication_mult_21_n24) );
  XOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U22 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_1__4_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_ab_0__5_), .Z(
        my_filter_adder_mult_8_multiplication_mult_21_n23) );
  XOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U21 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_1__5_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_ab_0__6_), .Z(
        my_filter_adder_mult_8_multiplication_mult_21_n22) );
  XOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U20 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_1__6_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_ab_0__7_), .Z(
        my_filter_adder_mult_8_multiplication_mult_21_n21) );
  XOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U19 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_1__7_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_ab_0__8_), .Z(
        my_filter_adder_mult_8_multiplication_mult_21_n20) );
  XOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U18 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_1__8_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_ab_0__9_), .Z(
        my_filter_adder_mult_8_multiplication_mult_21_n19) );
  XOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U17 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_1__9_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_ab_0__10_), .Z(
        my_filter_adder_mult_8_multiplication_mult_21_n18) );
  XOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U16 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_1__10_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_ab_0__11_), .Z(
        my_filter_adder_mult_8_multiplication_mult_21_n17) );
  XOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_U15 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_1__11_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_ab_0__12_), .Z(
        my_filter_adder_mult_8_multiplication_mult_21_n16) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S3_2_12 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_2__12_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_n15), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_ab_1__13_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_2__12_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_2__12_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_2_11 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_2__11_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_n4), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_n26), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_2__11_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_2__11_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_2_10 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_2__10_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_n5), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_n16), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_2__10_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_2__10_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_2_9 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_2__9_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_n6), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_n17), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_2__9_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_2__9_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_2_8 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_2__8_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_n7), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_n18), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_2__8_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_2__8_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_2_7 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_2__7_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_n8), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_n19), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_2__7_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_2__7_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_2_6 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_2__6_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_n9), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_n20), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_2__6_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_2__6_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_2_5 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_2__5_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_n10), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_n21), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_2__5_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_2__5_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_2_4 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_2__4_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_n11), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_n22), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_2__4_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_2__4_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_2_3 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_2__3_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_n12), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_n23), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_2__3_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_2__3_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_2_2 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_2__2_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_n13), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_n24), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_2__2_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_2__2_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_2_1 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_2__1_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_n14), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_n25), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_2__1_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_2__1_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S1_2_0 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_2__0_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_1__0_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_n27), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_2__0_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_A1_0_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S3_3_12 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_3__12_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_2__12_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_ab_2__13_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_3__12_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_3__12_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_3_11 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_3__11_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_2__11_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_2__12_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_3__11_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_3__11_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_3_10 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_3__10_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_2__10_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_2__11_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_3__10_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_3__10_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_3_9 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_3__9_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_2__9_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_2__10_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_3__9_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_3__9_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_3_8 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_3__8_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_2__8_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_2__9_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_3__8_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_3__8_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_3_7 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_3__7_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_2__7_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_2__8_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_3__7_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_3__7_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_3_6 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_3__6_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_2__6_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_2__7_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_3__6_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_3__6_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_3_5 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_3__5_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_2__5_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_2__6_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_3__5_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_3__5_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_3_4 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_3__4_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_2__4_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_2__5_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_3__4_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_3__4_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_3_3 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_3__3_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_2__3_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_2__4_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_3__3_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_3__3_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_3_2 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_3__2_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_2__2_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_2__3_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_3__2_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_3__2_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_3_1 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_3__1_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_2__1_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_2__2_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_3__1_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_3__1_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S1_3_0 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_3__0_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_2__0_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_2__1_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_3__0_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_A1_1_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S3_4_12 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_4__12_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_3__12_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_ab_3__13_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_4__12_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_4__12_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_4_11 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_4__11_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_3__11_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_3__12_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_4__11_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_4__11_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_4_10 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_4__10_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_3__10_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_3__11_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_4__10_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_4__10_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_4_9 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_4__9_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_3__9_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_3__10_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_4__9_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_4__9_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_4_8 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_4__8_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_3__8_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_3__9_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_4__8_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_4__8_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_4_7 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_4__7_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_3__7_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_3__8_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_4__7_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_4__7_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_4_6 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_4__6_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_3__6_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_3__7_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_4__6_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_4__6_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_4_5 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_4__5_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_3__5_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_3__6_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_4__5_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_4__5_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_4_4 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_4__4_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_3__4_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_3__5_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_4__4_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_4__4_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_4_3 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_4__3_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_3__3_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_3__4_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_4__3_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_4__3_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_4_2 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_4__2_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_3__2_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_3__3_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_4__2_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_4__2_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_4_1 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_4__1_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_3__1_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_3__2_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_4__1_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_4__1_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S1_4_0 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_4__0_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_3__0_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_3__1_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_4__0_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_A1_2_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S3_5_12 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_5__12_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_4__12_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_ab_4__13_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_5__12_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_5__12_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_5_11 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_5__11_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_4__11_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_4__12_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_5__11_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_5__11_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_5_10 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_5__10_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_4__10_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_4__11_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_5__10_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_5__10_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_5_9 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_5__9_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_4__9_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_4__10_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_5__9_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_5__9_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_5_8 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_5__8_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_4__8_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_4__9_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_5__8_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_5__8_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_5_7 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_5__7_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_4__7_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_4__8_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_5__7_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_5__7_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_5_6 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_5__6_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_4__6_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_4__7_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_5__6_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_5__6_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_5_5 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_5__5_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_4__5_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_4__6_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_5__5_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_5__5_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_5_4 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_5__4_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_4__4_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_4__5_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_5__4_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_5__4_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_5_3 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_5__3_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_4__3_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_4__4_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_5__3_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_5__3_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_5_2 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_5__2_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_4__2_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_4__3_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_5__2_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_5__2_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_5_1 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_5__1_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_4__1_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_4__2_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_5__1_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_5__1_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S1_5_0 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_5__0_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_4__0_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_4__1_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_5__0_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_A1_3_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S3_6_12 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_6__12_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_5__12_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_ab_5__13_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_6__12_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_6__12_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_6_11 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_6__11_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_5__11_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_5__12_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_6__11_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_6__11_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_6_10 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_6__10_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_5__10_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_5__11_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_6__10_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_6__10_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_6_9 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_6__9_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_5__9_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_5__10_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_6__9_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_6__9_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_6_8 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_6__8_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_5__8_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_5__9_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_6__8_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_6__8_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_6_7 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_6__7_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_5__7_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_5__8_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_6__7_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_6__7_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_6_6 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_6__6_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_5__6_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_5__7_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_6__6_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_6__6_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_6_5 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_6__5_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_5__5_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_5__6_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_6__5_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_6__5_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_6_4 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_6__4_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_5__4_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_5__5_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_6__4_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_6__4_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_6_3 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_6__3_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_5__3_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_5__4_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_6__3_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_6__3_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_6_2 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_6__2_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_5__2_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_5__3_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_6__2_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_6__2_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_6_1 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_6__1_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_5__1_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_5__2_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_6__1_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_6__1_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S1_6_0 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_6__0_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_5__0_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_5__1_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_6__0_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_A1_4_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S3_7_12 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_7__12_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_6__12_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_ab_6__13_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_7__12_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_7__12_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_7_11 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_7__11_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_6__11_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_6__12_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_7__11_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_7__11_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_7_10 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_7__10_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_6__10_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_6__11_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_7__10_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_7__10_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_7_9 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_7__9_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_6__9_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_6__10_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_7__9_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_7__9_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_7_8 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_7__8_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_6__8_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_6__9_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_7__8_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_7__8_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_7_7 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_7__7_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_6__7_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_6__8_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_7__7_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_7__7_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_7_6 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_7__6_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_6__6_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_6__7_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_7__6_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_7__6_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_7_5 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_7__5_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_6__5_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_6__6_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_7__5_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_7__5_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_7_4 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_7__4_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_6__4_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_6__5_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_7__4_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_7__4_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_7_3 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_7__3_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_6__3_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_6__4_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_7__3_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_7__3_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_7_2 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_7__2_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_6__2_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_6__3_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_7__2_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_7__2_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_7_1 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_7__1_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_6__1_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_6__2_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_7__1_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_7__1_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S1_7_0 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_7__0_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_6__0_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_6__1_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_7__0_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_A1_5_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S3_8_12 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_8__12_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_7__12_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_ab_7__13_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_8__12_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_8__12_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_8_11 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_8__11_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_7__11_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_7__12_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_8__11_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_8__11_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_8_10 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_8__10_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_7__10_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_7__11_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_8__10_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_8__10_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_8_9 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_8__9_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_7__9_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_7__10_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_8__9_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_8__9_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_8_8 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_8__8_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_7__8_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_7__9_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_8__8_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_8__8_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_8_7 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_8__7_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_7__7_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_7__8_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_8__7_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_8__7_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_8_6 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_8__6_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_7__6_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_7__7_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_8__6_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_8__6_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_8_5 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_8__5_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_7__5_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_7__6_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_8__5_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_8__5_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_8_4 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_8__4_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_7__4_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_7__5_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_8__4_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_8__4_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_8_3 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_8__3_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_7__3_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_7__4_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_8__3_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_8__3_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_8_2 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_8__2_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_7__2_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_7__3_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_8__2_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_8__2_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_8_1 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_8__1_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_7__1_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_7__2_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_8__1_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_8__1_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S1_8_0 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_8__0_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_7__0_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_7__1_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_8__0_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_A1_6_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S3_9_12 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_9__12_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_8__12_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_ab_8__13_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_9__12_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_9__12_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_9_11 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_9__11_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_8__11_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_8__12_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_9__11_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_9__11_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_9_10 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_9__10_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_8__10_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_8__11_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_9__10_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_9__10_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_9_9 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_9__9_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_8__9_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_8__10_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_9__9_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_9__9_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_9_8 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_9__8_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_8__8_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_8__9_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_9__8_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_9__8_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_9_7 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_9__7_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_8__7_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_8__8_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_9__7_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_9__7_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_9_6 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_9__6_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_8__6_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_8__7_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_9__6_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_9__6_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_9_5 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_9__5_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_8__5_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_8__6_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_9__5_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_9__5_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_9_4 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_9__4_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_8__4_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_8__5_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_9__4_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_9__4_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_9_3 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_9__3_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_8__3_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_8__4_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_9__3_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_9__3_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_9_2 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_9__2_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_8__2_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_8__3_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_9__2_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_9__2_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_9_1 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_9__1_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_8__1_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_8__2_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_9__1_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_9__1_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S1_9_0 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_9__0_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_8__0_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_8__1_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_9__0_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_A1_7_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S3_10_12 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_10__12_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_9__12_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_ab_9__13_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_10__12_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_10__12_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_10_11 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_10__11_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_9__11_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_9__12_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_10__11_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_10__11_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_10_10 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_10__10_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_9__10_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_9__11_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_10__10_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_10__10_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_10_9 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_10__9_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_9__9_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_9__10_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_10__9_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_10__9_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_10_8 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_10__8_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_9__8_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_9__9_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_10__8_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_10__8_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_10_7 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_10__7_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_9__7_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_9__8_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_10__7_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_10__7_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_10_6 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_10__6_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_9__6_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_9__7_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_10__6_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_10__6_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_10_5 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_10__5_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_9__5_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_9__6_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_10__5_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_10__5_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_10_4 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_10__4_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_9__4_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_9__5_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_10__4_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_10__4_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_10_3 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_10__3_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_9__3_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_9__4_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_10__3_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_10__3_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_10_2 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_10__2_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_9__2_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_9__3_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_10__2_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_10__2_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_10_1 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_10__1_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_9__1_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_9__2_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_10__1_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_10__1_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S1_10_0 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_10__0_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_9__0_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_9__1_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_10__0_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_A1_8_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S3_11_12 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_11__12_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_10__12_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_ab_10__13_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_11__12_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_11__12_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_11_11 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_11__11_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_10__11_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_10__12_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_11__11_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_11__11_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_11_10 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_11__10_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_10__10_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_10__11_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_11__10_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_11__10_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_11_9 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_11__9_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_10__9_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_10__10_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_11__9_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_11__9_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_11_8 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_11__8_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_10__8_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_10__9_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_11__8_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_11__8_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_11_7 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_11__7_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_10__7_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_10__8_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_11__7_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_11__7_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_11_6 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_11__6_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_10__6_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_10__7_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_11__6_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_11__6_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_11_5 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_11__5_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_10__5_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_10__6_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_11__5_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_11__5_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_11_4 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_11__4_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_10__4_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_10__5_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_11__4_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_11__4_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_11_3 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_11__3_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_10__3_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_10__4_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_11__3_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_11__3_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_11_2 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_11__2_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_10__2_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_10__3_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_11__2_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_11__2_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_11_1 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_11__1_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_10__1_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_10__2_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_11__1_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_11__1_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S1_11_0 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_11__0_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_10__0_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_10__1_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_11__0_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_A1_9_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S3_12_12 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_12__12_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_11__12_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_ab_11__13_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_12__12_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_12__12_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_12_11 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_12__11_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_11__11_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_11__12_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_12__11_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_12__11_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_12_10 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_12__10_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_11__10_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_11__11_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_12__10_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_12__10_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_12_9 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_12__9_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_11__9_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_11__10_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_12__9_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_12__9_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_12_8 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_12__8_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_11__8_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_11__9_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_12__8_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_12__8_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_12_7 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_12__7_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_11__7_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_11__8_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_12__7_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_12__7_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_12_6 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_12__6_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_11__6_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_11__7_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_12__6_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_12__6_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_12_5 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_12__5_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_11__5_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_11__6_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_12__5_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_12__5_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_12_4 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_12__4_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_11__4_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_11__5_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_12__4_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_12__4_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_12_3 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_12__3_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_11__3_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_11__4_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_12__3_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_12__3_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_12_2 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_12__2_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_11__2_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_11__3_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_12__2_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_12__2_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S2_12_1 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_12__1_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_11__1_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_11__2_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_12__1_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_12__1_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S1_12_0 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_12__0_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_11__0_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_11__1_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_12__0_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_A1_10_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S14_13 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_n86), .B(
        my_filter_adder_mult_8_multiplication_mult_21_n100), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_ab_13__13_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_13__13_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_13__13_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S5_12 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_13__12_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_12__12_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_ab_12__13_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_13__12_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_13__12_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S4_11 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_13__11_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_12__11_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_12__12_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_13__11_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_13__11_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S4_10 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_13__10_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_12__10_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_12__11_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_13__10_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_13__10_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S4_9 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_13__9_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_12__9_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_12__10_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_13__9_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_13__9_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S4_8 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_13__8_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_12__8_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_12__9_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_13__8_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_13__8_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S4_7 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_13__7_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_12__7_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_12__8_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_13__7_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_13__7_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S4_6 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_13__6_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_12__6_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_12__7_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_13__6_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_13__6_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S4_5 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_13__5_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_12__5_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_12__6_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_13__5_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_13__5_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S4_4 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_13__4_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_12__4_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_12__5_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_13__4_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_13__4_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S4_3 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_13__3_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_12__3_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_12__4_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_13__3_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_13__3_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S4_2 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_13__2_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_12__2_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_12__3_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_13__2_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_13__2_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S4_1 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_13__1_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_12__1_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_12__2_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_13__1_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_13__1_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S4_0 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_ab_13__0_), .B(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_12__0_), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_12__1_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_CARRYB_13__0_), .S(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_13__0_) );
  FA_X1 my_filter_adder_mult_8_multiplication_mult_21_S14_13_0 ( .A(
        my_filter_q_reg_chain_9__13_), .B(my_filter_q_reg_coeff[27]), .CI(
        my_filter_adder_mult_8_multiplication_mult_21_SUMB_13__0_), .CO(
        my_filter_adder_mult_8_multiplication_mult_21_A2_12_), .S(
        my_filter_adder_mult_8_res_mult[0]) );
  NAND2_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U72 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_A2_12_), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n28), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n56) );
  OAI21_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U71 ( .B1(
        my_filter_adder_mult_8_multiplication_mult_21_A2_12_), .B2(
        my_filter_adder_mult_8_multiplication_mult_21_n28), .A(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n56), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n59) );
  INV_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U70 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n59), .ZN(
        my_filter_adder_mult_8_res_mult[1]) );
  AND2_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U69 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n50), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n48), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n20) );
  AND2_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U68 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n49), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n43), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n28) );
  NAND2_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U66 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n47), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n44), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n17) );
  NAND2_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U65 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n46), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n42), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n25) );
  NAND2_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U64 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n45), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n41), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n33) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U63 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n47), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n44), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n15) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U61 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n46), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n42), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n23) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U60 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n45), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n41), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n31) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U59 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n50), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n48), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n21) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U58 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n49), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n43), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n29) );
  AND2_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U56 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n40), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n31), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n36) );
  AND2_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U55 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n35), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n30), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n44) );
  AND2_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U54 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n39), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n29), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n52) );
  NAND2_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U53 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n34), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n38), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n41) );
  NAND2_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U51 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n33), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n37), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n49) );
  NAND2_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U50 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n32), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n36), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n57) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U49 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n34), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n38), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n39) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U48 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n33), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n37), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n47) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U46 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n32), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n36), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n55) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U45 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n40), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n31), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n37) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U44 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n35), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n30), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n45) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U43 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_n39), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_n29), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n53) );
  OAI21_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U41 ( .B1(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n55), .B2(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n56), .A(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n57), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n51) );
  INV_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U40 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n55), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n60) );
  NAND2_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U39 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n60), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n57), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n58) );
  OAI21_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U38 ( .B1(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n15), .B2(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n16), .A(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n17), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n13) );
  OAI21_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U36 ( .B1(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n23), .B2(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n24), .A(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n25), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n19) );
  OAI21_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U35 ( .B1(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n31), .B2(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n32), .A(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n33), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n27) );
  OAI21_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U34 ( .B1(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n39), .B2(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n40), .A(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n41), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n35) );
  OAI21_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U33 ( .B1(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n47), .B2(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n48), .A(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n49), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n43) );
  INV_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U31 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n21), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n63) );
  AOI21_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U30 ( .B1(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n63), .B2(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n19), .A(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n20), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n16) );
  INV_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U29 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n29), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n71) );
  AOI21_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U28 ( .B1(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n71), .B2(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n27), .A(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n28), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n24) );
  INV_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U26 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n37), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n69) );
  AOI21_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U25 ( .B1(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n69), .B2(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n35), .A(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n36), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n32) );
  INV_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U24 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n45), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n67) );
  AOI21_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U23 ( .B1(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n67), .B2(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n43), .A(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n44), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n40) );
  INV_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U21 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n53), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n65) );
  AOI21_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U20 ( .B1(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n65), .B2(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n51), .A(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n52), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n48) );
  INV_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U19 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n15), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n62) );
  NAND2_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U18 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n62), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n17), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n18) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U16 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n20), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n21), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n22) );
  INV_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U13 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n23), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n64) );
  NAND2_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U12 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n64), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n25), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n26) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U11 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n28), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n29), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n30) );
  INV_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U10 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n31), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n70) );
  NAND2_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U9 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n70), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n33), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n34) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U8 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n36), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n37), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n38) );
  INV_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U7 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n39), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n68) );
  NAND2_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U6 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n68), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n41), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n42) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U5 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n44), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n45), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n46) );
  INV_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U4 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n47), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n66) );
  NAND2_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U3 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n66), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n49), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n50) );
  NOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U2 ( .A1(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n52), .A2(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n53), .ZN(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n54) );
  XOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U67 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n56), .B(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n58), .Z(
        my_filter_adder_mult_8_res_mult[2]) );
  XOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U62 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n51), .B(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n54), .Z(
        my_filter_adder_mult_8_res_mult[3]) );
  XOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U57 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n50), .B(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n48), .Z(
        my_filter_adder_mult_8_res_mult[4]) );
  XOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U52 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n43), .B(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n46), .Z(
        my_filter_adder_mult_8_res_mult[5]) );
  XOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U47 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n42), .B(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n40), .Z(
        my_filter_adder_mult_8_res_mult[6]) );
  XOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U42 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n35), .B(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n38), .Z(
        my_filter_adder_mult_8_res_mult[7]) );
  XOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U37 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n34), .B(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n32), .Z(
        my_filter_adder_mult_8_res_mult[8]) );
  XOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U32 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n27), .B(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n30), .Z(
        my_filter_adder_mult_8_res_mult[9]) );
  XOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U27 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n26), .B(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n24), .Z(
        my_filter_adder_mult_8_res_mult[10]) );
  XOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U22 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n19), .B(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n22), .Z(
        my_filter_adder_mult_8_res_mult[11]) );
  XOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U17 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n18), .B(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n16), .Z(
        my_filter_adder_mult_8_res_mult[12]) );
  XOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U15 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_n52), .B(
        my_filter_adder_mult_8_multiplication_mult_21_n51), .Z(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n14) );
  XOR2_X1 my_filter_adder_mult_8_multiplication_mult_21_FS_1_U14 ( .A(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n13), .B(
        my_filter_adder_mult_8_multiplication_mult_21_FS_1_n14), .Z(
        my_filter_adder_mult_8_res_mult[13]) );
  AND2_X1 my_filter_adder_mult_8_addition_add_19_U1 ( .A1(
        my_filter_data_sum[28]), .A2(my_filter_adder_mult_8_res_mult[0]), .ZN(
        my_filter_adder_mult_8_addition_add_19_n1) );
  XOR2_X1 my_filter_adder_mult_8_addition_add_19_U2 ( .A(
        my_filter_data_sum[28]), .B(my_filter_adder_mult_8_res_mult[0]), .Z(
        my_filter_data_sum[14]) );
  FA_X1 my_filter_adder_mult_8_addition_add_19_U1_1 ( .A(
        my_filter_adder_mult_8_res_mult[1]), .B(my_filter_data_sum[29]), .CI(
        my_filter_adder_mult_8_addition_add_19_n1), .CO(
        my_filter_adder_mult_8_addition_add_19_carry[2]), .S(
        my_filter_data_sum[15]) );
  FA_X1 my_filter_adder_mult_8_addition_add_19_U1_2 ( .A(
        my_filter_adder_mult_8_res_mult[2]), .B(my_filter_data_sum[30]), .CI(
        my_filter_adder_mult_8_addition_add_19_carry[2]), .CO(
        my_filter_adder_mult_8_addition_add_19_carry[3]), .S(
        my_filter_data_sum[16]) );
  FA_X1 my_filter_adder_mult_8_addition_add_19_U1_3 ( .A(
        my_filter_adder_mult_8_res_mult[3]), .B(my_filter_data_sum[31]), .CI(
        my_filter_adder_mult_8_addition_add_19_carry[3]), .CO(
        my_filter_adder_mult_8_addition_add_19_carry[4]), .S(
        my_filter_data_sum[17]) );
  FA_X1 my_filter_adder_mult_8_addition_add_19_U1_4 ( .A(
        my_filter_adder_mult_8_res_mult[4]), .B(my_filter_data_sum[32]), .CI(
        my_filter_adder_mult_8_addition_add_19_carry[4]), .CO(
        my_filter_adder_mult_8_addition_add_19_carry[5]), .S(
        my_filter_data_sum[18]) );
  FA_X1 my_filter_adder_mult_8_addition_add_19_U1_5 ( .A(
        my_filter_adder_mult_8_res_mult[5]), .B(my_filter_data_sum[33]), .CI(
        my_filter_adder_mult_8_addition_add_19_carry[5]), .CO(
        my_filter_adder_mult_8_addition_add_19_carry[6]), .S(
        my_filter_data_sum[19]) );
  FA_X1 my_filter_adder_mult_8_addition_add_19_U1_6 ( .A(
        my_filter_adder_mult_8_res_mult[6]), .B(my_filter_data_sum[34]), .CI(
        my_filter_adder_mult_8_addition_add_19_carry[6]), .CO(
        my_filter_adder_mult_8_addition_add_19_carry[7]), .S(
        my_filter_data_sum[20]) );
  FA_X1 my_filter_adder_mult_8_addition_add_19_U1_7 ( .A(
        my_filter_adder_mult_8_res_mult[7]), .B(my_filter_data_sum[35]), .CI(
        my_filter_adder_mult_8_addition_add_19_carry[7]), .CO(
        my_filter_adder_mult_8_addition_add_19_carry[8]), .S(
        my_filter_data_sum[21]) );
  FA_X1 my_filter_adder_mult_8_addition_add_19_U1_8 ( .A(
        my_filter_adder_mult_8_res_mult[8]), .B(my_filter_data_sum[36]), .CI(
        my_filter_adder_mult_8_addition_add_19_carry[8]), .CO(
        my_filter_adder_mult_8_addition_add_19_carry[9]), .S(
        my_filter_data_sum[22]) );
  FA_X1 my_filter_adder_mult_8_addition_add_19_U1_9 ( .A(
        my_filter_adder_mult_8_res_mult[9]), .B(my_filter_data_sum[37]), .CI(
        my_filter_adder_mult_8_addition_add_19_carry[9]), .CO(
        my_filter_adder_mult_8_addition_add_19_carry[10]), .S(
        my_filter_data_sum[23]) );
  FA_X1 my_filter_adder_mult_8_addition_add_19_U1_10 ( .A(
        my_filter_adder_mult_8_res_mult[10]), .B(my_filter_data_sum[38]), .CI(
        my_filter_adder_mult_8_addition_add_19_carry[10]), .CO(
        my_filter_adder_mult_8_addition_add_19_carry[11]), .S(
        my_filter_data_sum[24]) );
  FA_X1 my_filter_adder_mult_8_addition_add_19_U1_11 ( .A(
        my_filter_adder_mult_8_res_mult[11]), .B(my_filter_data_sum[39]), .CI(
        my_filter_adder_mult_8_addition_add_19_carry[11]), .CO(
        my_filter_adder_mult_8_addition_add_19_carry[12]), .S(
        my_filter_data_sum[25]) );
  FA_X1 my_filter_adder_mult_8_addition_add_19_U1_12 ( .A(
        my_filter_adder_mult_8_res_mult[12]), .B(my_filter_data_sum[40]), .CI(
        my_filter_adder_mult_8_addition_add_19_carry[12]), .CO(
        my_filter_adder_mult_8_addition_add_19_carry[13]), .S(
        my_filter_data_sum[26]) );
  FA_X1 my_filter_adder_mult_8_addition_add_19_U1_13 ( .A(
        my_filter_adder_mult_8_res_mult[13]), .B(my_filter_data_sum[41]), .CI(
        my_filter_adder_mult_8_addition_add_19_carry[13]), .S(
        my_filter_data_sum[27]) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U276 ( .A1(
        my_filter_q_reg_chain_10__11_), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_11__13_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U275 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_12__12_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U274 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_11__12_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U273 ( .A1(
        my_filter_q_reg_chain_10__10_), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_10__13_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U272 ( .A1(
        my_filter_q_reg_chain_10__9_), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_9__13_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U271 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_10__12_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U270 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n101), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_9__12_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U269 ( .A1(
        my_filter_q_reg_chain_10__8_), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_8__13_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U268 ( .A1(
        my_filter_q_reg_chain_10__7_), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_7__13_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U267 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_8__12_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U266 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_7__12_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U265 ( .A1(
        my_filter_q_reg_chain_10__6_), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_6__13_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U264 ( .A1(
        my_filter_q_reg_coeff[10]), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_13__10_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U263 ( .A1(
        my_filter_q_reg_coeff[11]), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_13__11_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U262 ( .A1(
        my_filter_q_reg_coeff[8]), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_13__8_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U261 ( .A1(
        my_filter_q_reg_coeff[9]), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_13__9_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U260 ( .A1(
        my_filter_q_reg_coeff[7]), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_13__7_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U259 ( .A1(
        my_filter_q_reg_coeff[12]), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_13__12_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U258 ( .A1(
        my_filter_q_reg_chain_10__12_), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_12__13_) );
  INV_X1 my_filter_adder_mult_9_multiplication_mult_21_U257 ( .A(
        my_filter_q_reg_chain_10__13_), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_n86) );
  INV_X1 my_filter_adder_mult_9_multiplication_mult_21_U256 ( .A(
        my_filter_q_reg_chain_10__9_), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_n90) );
  INV_X1 my_filter_adder_mult_9_multiplication_mult_21_U255 ( .A(
        my_filter_q_reg_chain_10__12_), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_n87) );
  INV_X1 my_filter_adder_mult_9_multiplication_mult_21_U254 ( .A(
        my_filter_q_reg_chain_10__11_), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_n88) );
  INV_X1 my_filter_adder_mult_9_multiplication_mult_21_U253 ( .A(
        my_filter_q_reg_chain_10__10_), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_n89) );
  INV_X1 my_filter_adder_mult_9_multiplication_mult_21_U252 ( .A(
        my_filter_q_reg_chain_10__8_), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_n91) );
  INV_X1 my_filter_adder_mult_9_multiplication_mult_21_U251 ( .A(
        my_filter_q_reg_chain_10__7_), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_n92) );
  INV_X1 my_filter_adder_mult_9_multiplication_mult_21_U250 ( .A(
        my_filter_q_reg_chain_10__6_), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_n93) );
  AND2_X1 my_filter_adder_mult_9_multiplication_mult_21_U249 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_ab_0__13_), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_ab_1__12_), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_n15) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U248 ( .A1(
        my_filter_q_reg_chain_10__1_), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_1__13_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U247 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_2__12_) );
  AND3_X1 my_filter_adder_mult_9_multiplication_mult_21_U246 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_ab_1__1_), .A2(
        my_filter_q_reg_coeff[0]), .A3(my_filter_q_reg_chain_10__0_), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_1__0_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U245 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_12__0_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U244 ( .A1(
        my_filter_q_reg_coeff[0]), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_13__0_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U243 ( .A1(
        my_filter_q_reg_chain_10__5_), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_5__13_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U242 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_6__12_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U241 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_5__12_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U240 ( .A1(
        my_filter_q_reg_chain_10__4_), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_4__13_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U239 ( .A1(
        my_filter_q_reg_chain_10__3_), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_3__13_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U238 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_4__12_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U237 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_3__12_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U236 ( .A1(
        my_filter_q_reg_chain_10__2_), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_2__13_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U235 ( .A1(
        my_filter_q_reg_coeff[6]), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_13__6_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U234 ( .A1(
        my_filter_q_reg_coeff[4]), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_13__4_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U233 ( .A1(
        my_filter_q_reg_coeff[5]), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_13__5_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U232 ( .A1(
        my_filter_q_reg_coeff[2]), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_13__2_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U231 ( .A1(
        my_filter_q_reg_coeff[3]), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_13__3_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U230 ( .A1(
        my_filter_q_reg_coeff[1]), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_13__1_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U229 ( .A1(
        my_filter_q_reg_chain_10__0_), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n100), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_0__13_) );
  INV_X1 my_filter_adder_mult_9_multiplication_mult_21_U228 ( .A(
        my_filter_q_reg_coeff[13]), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_n100) );
  INV_X1 my_filter_adder_mult_9_multiplication_mult_21_U227 ( .A(
        my_filter_q_reg_coeff[0]), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_n113) );
  INV_X1 my_filter_adder_mult_9_multiplication_mult_21_U226 ( .A(
        my_filter_q_reg_chain_10__0_), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_n99) );
  INV_X1 my_filter_adder_mult_9_multiplication_mult_21_U225 ( .A(
        my_filter_q_reg_coeff[1]), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_n112) );
  INV_X1 my_filter_adder_mult_9_multiplication_mult_21_U224 ( .A(
        my_filter_q_reg_chain_10__1_), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_n98) );
  INV_X1 my_filter_adder_mult_9_multiplication_mult_21_U223 ( .A(
        my_filter_q_reg_coeff[12]), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_n101) );
  INV_X1 my_filter_adder_mult_9_multiplication_mult_21_U222 ( .A(
        my_filter_q_reg_coeff[10]), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_n103) );
  INV_X1 my_filter_adder_mult_9_multiplication_mult_21_U221 ( .A(
        my_filter_q_reg_coeff[11]), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_n102) );
  INV_X1 my_filter_adder_mult_9_multiplication_mult_21_U220 ( .A(
        my_filter_q_reg_coeff[8]), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_n105) );
  INV_X1 my_filter_adder_mult_9_multiplication_mult_21_U219 ( .A(
        my_filter_q_reg_coeff[9]), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_n104) );
  INV_X1 my_filter_adder_mult_9_multiplication_mult_21_U218 ( .A(
        my_filter_q_reg_coeff[6]), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_n107) );
  INV_X1 my_filter_adder_mult_9_multiplication_mult_21_U217 ( .A(
        my_filter_q_reg_coeff[7]), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_n106) );
  INV_X1 my_filter_adder_mult_9_multiplication_mult_21_U216 ( .A(
        my_filter_q_reg_coeff[2]), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_n111) );
  INV_X1 my_filter_adder_mult_9_multiplication_mult_21_U215 ( .A(
        my_filter_q_reg_coeff[3]), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_n110) );
  INV_X1 my_filter_adder_mult_9_multiplication_mult_21_U214 ( .A(
        my_filter_q_reg_coeff[4]), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_n109) );
  INV_X1 my_filter_adder_mult_9_multiplication_mult_21_U213 ( .A(
        my_filter_q_reg_coeff[5]), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_n108) );
  INV_X1 my_filter_adder_mult_9_multiplication_mult_21_U212 ( .A(
        my_filter_q_reg_chain_10__5_), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_n94) );
  INV_X1 my_filter_adder_mult_9_multiplication_mult_21_U211 ( .A(
        my_filter_q_reg_chain_10__4_), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_n95) );
  INV_X1 my_filter_adder_mult_9_multiplication_mult_21_U210 ( .A(
        my_filter_q_reg_chain_10__3_), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_n96) );
  INV_X1 my_filter_adder_mult_9_multiplication_mult_21_U209 ( .A(
        my_filter_q_reg_chain_10__2_), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_n97) );
  AND2_X1 my_filter_adder_mult_9_multiplication_mult_21_U208 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_13__12_), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_13__13_), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_n3) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U207 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n100), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n86), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_13__13_) );
  AND2_X1 my_filter_adder_mult_9_multiplication_mult_21_U206 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_13__9_), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_13__10_), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_n52) );
  AND2_X1 my_filter_adder_mult_9_multiplication_mult_21_U205 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_13__7_), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_13__8_), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_n51) );
  AND2_X1 my_filter_adder_mult_9_multiplication_mult_21_U204 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_13__5_), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_13__6_), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_n50) );
  AND2_X1 my_filter_adder_mult_9_multiplication_mult_21_U203 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_13__10_), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_13__11_), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_n48) );
  AND2_X1 my_filter_adder_mult_9_multiplication_mult_21_U202 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_13__8_), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_13__9_), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_n47) );
  AND2_X1 my_filter_adder_mult_9_multiplication_mult_21_U201 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_13__6_), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_13__7_), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_n46) );
  AND2_X1 my_filter_adder_mult_9_multiplication_mult_21_U200 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_13__4_), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_13__5_), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_n37) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U199 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_12__11_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U198 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_12__9_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U197 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_12__10_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U196 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_11__10_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U195 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_11__11_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U194 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_10__11_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U193 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_12__8_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U192 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_11__9_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U191 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_10__10_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U190 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n102), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_9__11_) );
  AND2_X1 my_filter_adder_mult_9_multiplication_mult_21_U189 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_13__11_), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_13__12_), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_n27) );
  AND2_X1 my_filter_adder_mult_9_multiplication_mult_21_U188 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_13__3_), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_13__4_), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_n38) );
  AND2_X1 my_filter_adder_mult_9_multiplication_mult_21_U187 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_13__1_), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_13__2_), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_n39) );
  AND2_X1 my_filter_adder_mult_9_multiplication_mult_21_U186 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_13__2_), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_13__3_), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_n36) );
  AND2_X1 my_filter_adder_mult_9_multiplication_mult_21_U185 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_13__0_), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_13__1_), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_n35) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U184 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_12__1_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U183 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_10__0_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U182 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_11__0_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U181 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_11__1_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U180 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_10__1_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U179 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_8__0_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U178 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n113), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_9__0_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U177 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n112), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_9__1_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U176 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n110), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_9__3_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U175 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_8__1_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U174 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_8__3_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U173 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_6__0_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U172 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_7__0_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U171 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_7__1_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U170 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_7__3_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U169 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_7__5_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U168 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_6__1_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U167 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_6__3_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U166 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_6__5_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U165 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_4__0_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U164 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_5__0_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U163 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_5__1_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U162 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_5__3_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U161 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_5__5_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U160 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_5__7_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U159 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_4__1_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U158 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_4__3_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U157 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_4__5_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U156 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_4__7_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U155 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_2__0_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U154 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n113), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_3__0_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U153 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_3__1_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U152 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_3__3_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U151 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_3__5_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U150 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_3__7_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U149 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_3__9_) );
  AND2_X1 my_filter_adder_mult_9_multiplication_mult_21_U148 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_ab_0__2_), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_ab_1__1_), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_n14) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U147 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n112), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_2__1_) );
  AND2_X1 my_filter_adder_mult_9_multiplication_mult_21_U146 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_ab_0__4_), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_ab_1__3_), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_n12) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U145 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_2__3_) );
  AND2_X1 my_filter_adder_mult_9_multiplication_mult_21_U144 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_ab_0__6_), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_ab_1__5_), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_n10) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U143 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_2__5_) );
  AND2_X1 my_filter_adder_mult_9_multiplication_mult_21_U142 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_ab_0__8_), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_ab_1__7_), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_n8) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U141 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_2__7_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U140 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_12__7_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U139 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_11__8_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U138 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_10__9_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U137 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_12__5_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U136 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_12__6_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U135 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n103), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_9__10_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U134 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_11__6_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U133 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_11__7_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U132 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_8__11_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U131 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_10__7_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U130 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_10__8_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U129 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_12__3_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U128 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_12__4_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U127 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n105), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_9__8_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U126 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n104), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_9__9_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U125 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_11__4_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U124 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_11__5_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U123 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n87), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_12__2_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U122 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_8__9_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U121 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_8__10_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U120 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_10__5_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U119 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_10__6_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U118 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_11__3_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U117 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_7__10_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U116 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_7__11_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U115 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n107), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_9__6_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U114 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n106), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_9__7_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U113 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n88), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_11__2_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U112 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_10__4_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U111 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_6__11_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U110 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_8__7_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U109 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_8__8_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U108 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_10__2_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U107 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n89), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_10__3_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U106 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n108), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_9__5_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U105 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_7__8_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U104 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_7__9_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U103 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n111), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_9__2_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U102 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n90), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n109), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_9__4_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U101 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_8__6_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U100 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_6__9_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U99 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_6__10_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U98 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_8__2_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U97 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_8__4_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U96 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n91), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_8__5_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U95 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_7__7_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U94 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_5__10_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U93 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_5__11_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U92 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_7__2_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U91 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_7__4_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U90 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n92), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_7__6_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U89 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_6__8_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U88 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_4__11_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U87 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_6__2_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U86 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_6__4_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U85 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_6__6_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U84 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n93), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_6__7_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U83 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_5__9_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U82 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_5__2_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U81 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_5__4_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U80 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_5__6_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U79 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n94), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_5__8_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U78 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_4__10_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U77 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_4__2_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U76 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_4__4_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U75 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_4__6_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U74 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_4__8_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U73 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n95), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_4__9_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U72 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_3__11_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U71 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_3__2_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U70 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_3__4_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U69 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_3__6_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U68 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_3__8_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U67 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n96), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_3__10_) );
  AND2_X1 my_filter_adder_mult_9_multiplication_mult_21_U66 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_ab_0__3_), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_ab_1__2_), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_n13) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U65 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_2__2_) );
  AND2_X1 my_filter_adder_mult_9_multiplication_mult_21_U64 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_ab_0__5_), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_ab_1__4_), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_n11) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U63 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_2__4_) );
  AND2_X1 my_filter_adder_mult_9_multiplication_mult_21_U62 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_ab_0__7_), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_ab_1__6_), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_n9) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U61 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_2__6_) );
  AND2_X1 my_filter_adder_mult_9_multiplication_mult_21_U60 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_ab_0__9_), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_ab_1__8_), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_n7) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U59 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_2__8_) );
  AND2_X1 my_filter_adder_mult_9_multiplication_mult_21_U58 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_ab_0__10_), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_ab_1__9_), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_n6) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U57 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_2__9_) );
  AND2_X1 my_filter_adder_mult_9_multiplication_mult_21_U56 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_ab_0__11_), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_ab_1__10_), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_n5) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U55 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_2__10_) );
  AND2_X1 my_filter_adder_mult_9_multiplication_mult_21_U54 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_ab_0__12_), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_ab_1__11_), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_n4) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U52 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n97), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_2__11_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U51 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_1__12_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U50 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_1__2_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U48 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_1__3_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U47 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_1__4_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U46 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_1__5_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U39 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_1__6_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U38 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_1__7_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U37 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_1__8_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U36 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_1__9_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U35 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_1__10_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U26 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n98), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_1__11_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U14 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n111), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_0__2_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U13 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n110), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_0__3_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U12 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n109), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_0__4_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U11 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n108), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_0__5_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U10 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n107), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_0__6_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U9 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n106), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_0__7_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U8 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n105), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_0__8_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U7 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n104), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_0__9_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U6 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n103), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_0__10_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U5 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n102), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_0__11_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U4 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n101), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n99), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_0__12_) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U3 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n98), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n112), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_ab_1__1_) );
  INV_X1 my_filter_adder_mult_9_multiplication_mult_21_U2 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_13__13_), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_n85) );
  XOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U49 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_13__10_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_13__11_), .Z(
        my_filter_adder_mult_9_multiplication_mult_21_n49) );
  XOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U45 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_13__11_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_13__12_), .Z(
        my_filter_adder_mult_9_multiplication_mult_21_n45) );
  XOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U44 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_13__8_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_13__9_), .Z(
        my_filter_adder_mult_9_multiplication_mult_21_n44) );
  XOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U43 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_13__9_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_13__10_), .Z(
        my_filter_adder_mult_9_multiplication_mult_21_n43) );
  XOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U42 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_13__6_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_13__7_), .Z(
        my_filter_adder_mult_9_multiplication_mult_21_n42) );
  XOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U41 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_13__7_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_13__8_), .Z(
        my_filter_adder_mult_9_multiplication_mult_21_n41) );
  XOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U40 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_13__12_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_13__13_), .Z(
        my_filter_adder_mult_9_multiplication_mult_21_n40) );
  XOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U34 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_13__4_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_13__5_), .Z(
        my_filter_adder_mult_9_multiplication_mult_21_n34) );
  XOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U33 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_13__5_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_13__6_), .Z(
        my_filter_adder_mult_9_multiplication_mult_21_n33) );
  XOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U32 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_13__2_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_13__3_), .Z(
        my_filter_adder_mult_9_multiplication_mult_21_n32) );
  XOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U31 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_13__3_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_13__4_), .Z(
        my_filter_adder_mult_9_multiplication_mult_21_n31) );
  XOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U30 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_13__0_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_13__1_), .Z(
        my_filter_adder_mult_9_multiplication_mult_21_n30) );
  XOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U29 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_13__1_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_13__2_), .Z(
        my_filter_adder_mult_9_multiplication_mult_21_n29) );
  XOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U27 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_1__1_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_ab_0__2_), .Z(
        my_filter_adder_mult_9_multiplication_mult_21_n28) );
  XOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U25 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_1__12_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_ab_0__13_), .Z(
        my_filter_adder_mult_9_multiplication_mult_21_n26) );
  XOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U24 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_1__2_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_ab_0__3_), .Z(
        my_filter_adder_mult_9_multiplication_mult_21_n25) );
  XOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U23 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_1__3_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_ab_0__4_), .Z(
        my_filter_adder_mult_9_multiplication_mult_21_n24) );
  XOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U22 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_1__4_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_ab_0__5_), .Z(
        my_filter_adder_mult_9_multiplication_mult_21_n23) );
  XOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U21 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_1__5_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_ab_0__6_), .Z(
        my_filter_adder_mult_9_multiplication_mult_21_n22) );
  XOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U20 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_1__6_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_ab_0__7_), .Z(
        my_filter_adder_mult_9_multiplication_mult_21_n21) );
  XOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U19 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_1__7_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_ab_0__8_), .Z(
        my_filter_adder_mult_9_multiplication_mult_21_n20) );
  XOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U18 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_1__8_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_ab_0__9_), .Z(
        my_filter_adder_mult_9_multiplication_mult_21_n19) );
  XOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U17 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_1__9_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_ab_0__10_), .Z(
        my_filter_adder_mult_9_multiplication_mult_21_n18) );
  XOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U16 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_1__10_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_ab_0__11_), .Z(
        my_filter_adder_mult_9_multiplication_mult_21_n17) );
  XOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_U15 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_1__11_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_ab_0__12_), .Z(
        my_filter_adder_mult_9_multiplication_mult_21_n16) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S3_2_12 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_2__12_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_n15), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_ab_1__13_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_2__12_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_2__12_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_2_11 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_2__11_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_n4), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_n26), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_2__11_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_2__11_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_2_10 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_2__10_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_n5), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_n16), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_2__10_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_2__10_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_2_9 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_2__9_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_n6), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_n17), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_2__9_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_2__9_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_2_8 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_2__8_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_n7), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_n18), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_2__8_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_2__8_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_2_7 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_2__7_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_n8), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_n19), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_2__7_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_2__7_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_2_6 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_2__6_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_n9), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_n20), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_2__6_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_2__6_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_2_5 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_2__5_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_n10), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_n21), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_2__5_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_2__5_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_2_4 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_2__4_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_n11), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_n22), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_2__4_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_2__4_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_2_3 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_2__3_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_n12), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_n23), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_2__3_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_2__3_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_2_2 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_2__2_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_n13), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_n24), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_2__2_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_2__2_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_2_1 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_2__1_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_n14), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_n25), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_2__1_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_2__1_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S1_2_0 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_2__0_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_1__0_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_n28), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_2__0_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_A1_0_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S3_3_12 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_3__12_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_2__12_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_ab_2__13_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_3__12_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_3__12_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_3_11 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_3__11_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_2__11_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_2__12_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_3__11_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_3__11_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_3_10 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_3__10_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_2__10_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_2__11_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_3__10_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_3__10_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_3_9 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_3__9_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_2__9_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_2__10_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_3__9_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_3__9_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_3_8 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_3__8_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_2__8_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_2__9_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_3__8_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_3__8_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_3_7 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_3__7_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_2__7_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_2__8_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_3__7_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_3__7_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_3_6 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_3__6_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_2__6_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_2__7_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_3__6_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_3__6_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_3_5 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_3__5_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_2__5_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_2__6_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_3__5_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_3__5_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_3_4 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_3__4_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_2__4_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_2__5_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_3__4_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_3__4_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_3_3 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_3__3_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_2__3_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_2__4_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_3__3_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_3__3_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_3_2 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_3__2_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_2__2_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_2__3_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_3__2_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_3__2_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_3_1 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_3__1_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_2__1_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_2__2_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_3__1_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_3__1_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S1_3_0 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_3__0_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_2__0_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_2__1_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_3__0_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_A1_1_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S3_4_12 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_4__12_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_3__12_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_ab_3__13_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_4__12_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_4__12_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_4_11 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_4__11_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_3__11_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_3__12_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_4__11_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_4__11_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_4_10 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_4__10_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_3__10_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_3__11_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_4__10_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_4__10_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_4_9 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_4__9_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_3__9_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_3__10_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_4__9_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_4__9_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_4_8 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_4__8_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_3__8_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_3__9_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_4__8_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_4__8_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_4_7 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_4__7_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_3__7_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_3__8_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_4__7_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_4__7_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_4_6 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_4__6_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_3__6_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_3__7_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_4__6_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_4__6_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_4_5 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_4__5_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_3__5_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_3__6_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_4__5_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_4__5_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_4_4 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_4__4_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_3__4_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_3__5_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_4__4_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_4__4_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_4_3 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_4__3_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_3__3_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_3__4_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_4__3_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_4__3_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_4_2 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_4__2_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_3__2_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_3__3_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_4__2_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_4__2_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_4_1 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_4__1_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_3__1_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_3__2_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_4__1_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_4__1_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S1_4_0 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_4__0_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_3__0_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_3__1_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_4__0_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_A1_2_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S3_5_12 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_5__12_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_4__12_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_ab_4__13_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_5__12_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_5__12_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_5_11 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_5__11_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_4__11_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_4__12_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_5__11_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_5__11_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_5_10 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_5__10_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_4__10_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_4__11_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_5__10_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_5__10_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_5_9 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_5__9_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_4__9_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_4__10_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_5__9_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_5__9_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_5_8 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_5__8_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_4__8_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_4__9_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_5__8_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_5__8_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_5_7 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_5__7_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_4__7_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_4__8_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_5__7_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_5__7_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_5_6 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_5__6_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_4__6_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_4__7_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_5__6_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_5__6_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_5_5 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_5__5_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_4__5_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_4__6_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_5__5_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_5__5_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_5_4 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_5__4_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_4__4_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_4__5_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_5__4_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_5__4_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_5_3 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_5__3_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_4__3_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_4__4_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_5__3_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_5__3_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_5_2 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_5__2_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_4__2_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_4__3_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_5__2_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_5__2_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_5_1 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_5__1_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_4__1_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_4__2_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_5__1_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_5__1_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S1_5_0 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_5__0_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_4__0_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_4__1_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_5__0_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_A1_3_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S3_6_12 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_6__12_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_5__12_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_ab_5__13_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_6__12_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_6__12_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_6_11 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_6__11_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_5__11_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_5__12_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_6__11_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_6__11_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_6_10 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_6__10_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_5__10_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_5__11_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_6__10_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_6__10_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_6_9 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_6__9_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_5__9_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_5__10_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_6__9_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_6__9_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_6_8 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_6__8_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_5__8_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_5__9_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_6__8_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_6__8_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_6_7 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_6__7_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_5__7_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_5__8_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_6__7_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_6__7_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_6_6 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_6__6_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_5__6_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_5__7_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_6__6_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_6__6_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_6_5 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_6__5_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_5__5_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_5__6_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_6__5_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_6__5_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_6_4 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_6__4_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_5__4_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_5__5_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_6__4_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_6__4_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_6_3 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_6__3_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_5__3_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_5__4_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_6__3_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_6__3_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_6_2 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_6__2_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_5__2_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_5__3_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_6__2_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_6__2_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_6_1 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_6__1_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_5__1_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_5__2_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_6__1_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_6__1_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S1_6_0 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_6__0_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_5__0_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_5__1_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_6__0_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_A1_4_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S3_7_12 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_7__12_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_6__12_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_ab_6__13_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_7__12_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_7__12_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_7_11 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_7__11_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_6__11_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_6__12_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_7__11_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_7__11_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_7_10 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_7__10_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_6__10_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_6__11_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_7__10_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_7__10_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_7_9 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_7__9_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_6__9_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_6__10_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_7__9_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_7__9_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_7_8 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_7__8_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_6__8_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_6__9_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_7__8_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_7__8_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_7_7 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_7__7_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_6__7_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_6__8_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_7__7_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_7__7_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_7_6 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_7__6_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_6__6_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_6__7_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_7__6_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_7__6_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_7_5 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_7__5_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_6__5_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_6__6_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_7__5_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_7__5_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_7_4 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_7__4_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_6__4_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_6__5_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_7__4_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_7__4_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_7_3 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_7__3_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_6__3_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_6__4_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_7__3_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_7__3_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_7_2 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_7__2_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_6__2_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_6__3_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_7__2_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_7__2_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_7_1 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_7__1_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_6__1_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_6__2_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_7__1_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_7__1_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S1_7_0 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_7__0_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_6__0_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_6__1_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_7__0_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_A1_5_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S3_8_12 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_8__12_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_7__12_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_ab_7__13_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_8__12_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_8__12_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_8_11 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_8__11_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_7__11_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_7__12_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_8__11_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_8__11_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_8_10 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_8__10_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_7__10_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_7__11_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_8__10_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_8__10_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_8_9 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_8__9_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_7__9_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_7__10_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_8__9_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_8__9_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_8_8 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_8__8_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_7__8_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_7__9_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_8__8_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_8__8_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_8_7 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_8__7_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_7__7_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_7__8_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_8__7_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_8__7_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_8_6 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_8__6_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_7__6_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_7__7_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_8__6_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_8__6_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_8_5 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_8__5_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_7__5_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_7__6_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_8__5_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_8__5_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_8_4 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_8__4_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_7__4_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_7__5_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_8__4_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_8__4_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_8_3 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_8__3_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_7__3_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_7__4_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_8__3_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_8__3_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_8_2 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_8__2_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_7__2_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_7__3_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_8__2_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_8__2_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_8_1 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_8__1_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_7__1_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_7__2_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_8__1_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_8__1_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S1_8_0 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_8__0_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_7__0_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_7__1_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_8__0_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_A1_6_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S3_9_12 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_9__12_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_8__12_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_ab_8__13_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_9__12_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_9__12_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_9_11 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_9__11_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_8__11_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_8__12_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_9__11_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_9__11_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_9_10 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_9__10_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_8__10_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_8__11_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_9__10_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_9__10_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_9_9 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_9__9_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_8__9_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_8__10_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_9__9_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_9__9_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_9_8 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_9__8_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_8__8_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_8__9_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_9__8_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_9__8_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_9_7 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_9__7_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_8__7_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_8__8_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_9__7_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_9__7_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_9_6 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_9__6_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_8__6_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_8__7_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_9__6_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_9__6_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_9_5 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_9__5_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_8__5_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_8__6_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_9__5_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_9__5_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_9_4 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_9__4_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_8__4_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_8__5_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_9__4_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_9__4_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_9_3 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_9__3_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_8__3_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_8__4_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_9__3_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_9__3_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_9_2 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_9__2_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_8__2_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_8__3_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_9__2_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_9__2_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_9_1 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_9__1_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_8__1_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_8__2_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_9__1_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_9__1_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S1_9_0 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_9__0_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_8__0_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_8__1_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_9__0_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_A1_7_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S3_10_12 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_10__12_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_9__12_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_ab_9__13_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_10__12_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_10__12_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_10_11 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_10__11_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_9__11_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_9__12_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_10__11_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_10__11_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_10_10 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_10__10_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_9__10_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_9__11_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_10__10_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_10__10_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_10_9 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_10__9_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_9__9_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_9__10_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_10__9_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_10__9_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_10_8 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_10__8_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_9__8_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_9__9_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_10__8_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_10__8_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_10_7 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_10__7_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_9__7_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_9__8_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_10__7_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_10__7_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_10_6 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_10__6_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_9__6_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_9__7_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_10__6_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_10__6_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_10_5 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_10__5_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_9__5_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_9__6_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_10__5_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_10__5_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_10_4 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_10__4_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_9__4_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_9__5_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_10__4_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_10__4_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_10_3 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_10__3_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_9__3_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_9__4_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_10__3_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_10__3_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_10_2 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_10__2_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_9__2_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_9__3_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_10__2_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_10__2_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_10_1 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_10__1_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_9__1_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_9__2_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_10__1_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_10__1_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S1_10_0 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_10__0_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_9__0_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_9__1_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_10__0_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_A1_8_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S3_11_12 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_11__12_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_10__12_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_ab_10__13_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_11__12_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_11__12_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_11_11 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_11__11_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_10__11_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_10__12_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_11__11_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_11__11_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_11_10 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_11__10_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_10__10_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_10__11_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_11__10_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_11__10_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_11_9 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_11__9_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_10__9_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_10__10_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_11__9_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_11__9_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_11_8 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_11__8_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_10__8_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_10__9_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_11__8_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_11__8_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_11_7 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_11__7_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_10__7_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_10__8_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_11__7_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_11__7_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_11_6 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_11__6_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_10__6_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_10__7_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_11__6_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_11__6_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_11_5 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_11__5_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_10__5_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_10__6_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_11__5_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_11__5_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_11_4 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_11__4_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_10__4_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_10__5_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_11__4_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_11__4_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_11_3 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_11__3_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_10__3_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_10__4_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_11__3_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_11__3_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_11_2 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_11__2_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_10__2_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_10__3_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_11__2_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_11__2_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_11_1 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_11__1_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_10__1_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_10__2_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_11__1_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_11__1_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S1_11_0 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_11__0_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_10__0_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_10__1_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_11__0_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_A1_9_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S3_12_12 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_12__12_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_11__12_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_ab_11__13_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_12__12_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_12__12_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_12_11 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_12__11_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_11__11_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_11__12_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_12__11_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_12__11_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_12_10 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_12__10_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_11__10_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_11__11_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_12__10_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_12__10_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_12_9 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_12__9_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_11__9_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_11__10_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_12__9_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_12__9_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_12_8 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_12__8_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_11__8_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_11__9_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_12__8_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_12__8_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_12_7 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_12__7_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_11__7_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_11__8_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_12__7_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_12__7_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_12_6 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_12__6_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_11__6_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_11__7_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_12__6_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_12__6_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_12_5 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_12__5_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_11__5_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_11__6_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_12__5_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_12__5_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_12_4 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_12__4_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_11__4_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_11__5_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_12__4_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_12__4_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_12_3 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_12__3_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_11__3_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_11__4_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_12__3_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_12__3_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_12_2 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_12__2_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_11__2_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_11__3_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_12__2_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_12__2_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S2_12_1 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_12__1_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_11__1_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_11__2_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_12__1_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_12__1_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S1_12_0 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_12__0_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_11__0_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_11__1_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_12__0_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_A1_10_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S14_13 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_n86), .B(
        my_filter_adder_mult_9_multiplication_mult_21_n100), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_ab_13__13_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_13__13_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_13__13_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S5_12 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_13__12_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_12__12_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_ab_12__13_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_13__12_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_13__12_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S4_11 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_13__11_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_12__11_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_12__12_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_13__11_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_13__11_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S4_10 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_13__10_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_12__10_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_12__11_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_13__10_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_13__10_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S4_9 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_13__9_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_12__9_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_12__10_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_13__9_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_13__9_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S4_8 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_13__8_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_12__8_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_12__9_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_13__8_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_13__8_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S4_7 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_13__7_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_12__7_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_12__8_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_13__7_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_13__7_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S4_6 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_13__6_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_12__6_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_12__7_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_13__6_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_13__6_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S4_5 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_13__5_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_12__5_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_12__6_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_13__5_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_13__5_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S4_4 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_13__4_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_12__4_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_12__5_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_13__4_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_13__4_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S4_3 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_13__3_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_12__3_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_12__4_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_13__3_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_13__3_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S4_2 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_13__2_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_12__2_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_12__3_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_13__2_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_13__2_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S4_1 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_13__1_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_12__1_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_12__2_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_13__1_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_13__1_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S4_0 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_ab_13__0_), .B(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_12__0_), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_12__1_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_CARRYB_13__0_), .S(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_13__0_) );
  FA_X1 my_filter_adder_mult_9_multiplication_mult_21_S14_13_0 ( .A(
        my_filter_q_reg_chain_10__13_), .B(my_filter_q_reg_coeff[13]), .CI(
        my_filter_adder_mult_9_multiplication_mult_21_SUMB_13__0_), .CO(
        my_filter_adder_mult_9_multiplication_mult_21_A2_12_), .S(
        my_filter_adder_mult_9_res_mult[0]) );
  NAND2_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U72 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_A2_12_), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n30), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n56) );
  OAI21_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U71 ( .B1(
        my_filter_adder_mult_9_multiplication_mult_21_A2_12_), .B2(
        my_filter_adder_mult_9_multiplication_mult_21_n30), .A(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n56), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n59) );
  INV_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U70 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n59), .ZN(
        my_filter_adder_mult_9_res_mult[1]) );
  AND2_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U69 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n52), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n49), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n20) );
  AND2_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U68 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n51), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n44), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n28) );
  AND2_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U66 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n50), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n42), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n36) );
  NAND2_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U65 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n48), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n45), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n17) );
  NAND2_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U64 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n47), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n43), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n25) );
  NAND2_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U63 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n46), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n41), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n33) );
  NAND2_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U61 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n37), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n33), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n41) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U60 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n48), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n45), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n15) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U59 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n47), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n43), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n23) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U58 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n46), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n41), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n31) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U56 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n52), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n49), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n21) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U55 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n51), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n44), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n29) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U54 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n50), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n42), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n37) );
  AND2_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U53 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n38), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n34), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n44) );
  AND2_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U51 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n39), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n32), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n52) );
  NAND2_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U50 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n36), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n31), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n49) );
  NAND2_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U49 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n35), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n29), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n57) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U48 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n37), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n33), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n39) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U46 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n36), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n31), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n47) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U45 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n35), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n29), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n55) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U44 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n38), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n34), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n45) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U43 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_n39), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_n32), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n53) );
  OAI21_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U41 ( .B1(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n55), .B2(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n56), .A(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n57), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n51) );
  INV_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U40 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n55), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n60) );
  NAND2_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U39 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n60), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n57), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n58) );
  OAI21_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U38 ( .B1(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n15), .B2(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n16), .A(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n17), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n13) );
  OAI21_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U36 ( .B1(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n23), .B2(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n24), .A(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n25), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n19) );
  OAI21_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U35 ( .B1(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n31), .B2(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n32), .A(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n33), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n27) );
  OAI21_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U34 ( .B1(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n39), .B2(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n40), .A(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n41), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n35) );
  OAI21_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U33 ( .B1(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n47), .B2(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n48), .A(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n49), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n43) );
  INV_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U31 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n21), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n63) );
  AOI21_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U30 ( .B1(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n63), .B2(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n19), .A(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n20), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n16) );
  INV_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U29 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n29), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n71) );
  AOI21_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U28 ( .B1(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n71), .B2(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n27), .A(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n28), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n24) );
  INV_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U26 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n37), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n69) );
  AOI21_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U25 ( .B1(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n69), .B2(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n35), .A(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n36), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n32) );
  INV_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U24 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n45), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n67) );
  AOI21_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U23 ( .B1(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n67), .B2(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n43), .A(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n44), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n40) );
  INV_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U21 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n53), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n65) );
  AOI21_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U20 ( .B1(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n65), .B2(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n51), .A(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n52), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n48) );
  INV_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U19 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n15), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n62) );
  NAND2_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U18 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n62), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n17), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n18) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U16 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n20), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n21), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n22) );
  INV_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U13 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n23), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n64) );
  NAND2_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U12 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n64), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n25), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n26) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U11 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n28), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n29), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n30) );
  INV_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U10 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n31), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n70) );
  NAND2_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U9 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n70), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n33), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n34) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U8 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n36), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n37), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n38) );
  INV_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U7 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n39), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n68) );
  NAND2_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U6 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n68), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n41), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n42) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U5 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n44), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n45), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n46) );
  INV_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U4 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n47), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n66) );
  NAND2_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U3 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n66), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n49), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n50) );
  NOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U2 ( .A1(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n52), .A2(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n53), .ZN(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n54) );
  XOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U67 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n56), .B(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n58), .Z(
        my_filter_adder_mult_9_res_mult[2]) );
  XOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U62 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n51), .B(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n54), .Z(
        my_filter_adder_mult_9_res_mult[3]) );
  XOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U57 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n50), .B(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n48), .Z(
        my_filter_adder_mult_9_res_mult[4]) );
  XOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U52 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n43), .B(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n46), .Z(
        my_filter_adder_mult_9_res_mult[5]) );
  XOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U47 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n42), .B(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n40), .Z(
        my_filter_adder_mult_9_res_mult[6]) );
  XOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U42 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n35), .B(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n38), .Z(
        my_filter_adder_mult_9_res_mult[7]) );
  XOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U37 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n34), .B(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n32), .Z(
        my_filter_adder_mult_9_res_mult[8]) );
  XOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U32 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n27), .B(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n30), .Z(
        my_filter_adder_mult_9_res_mult[9]) );
  XOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U27 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n26), .B(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n24), .Z(
        my_filter_adder_mult_9_res_mult[10]) );
  XOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U22 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n19), .B(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n22), .Z(
        my_filter_adder_mult_9_res_mult[11]) );
  XOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U17 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n18), .B(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n16), .Z(
        my_filter_adder_mult_9_res_mult[12]) );
  XOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U15 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_n27), .B(
        my_filter_adder_mult_9_multiplication_mult_21_n40), .Z(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n14) );
  XOR2_X1 my_filter_adder_mult_9_multiplication_mult_21_FS_1_U14 ( .A(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n13), .B(
        my_filter_adder_mult_9_multiplication_mult_21_FS_1_n14), .Z(
        my_filter_adder_mult_9_res_mult[13]) );
  AND2_X1 my_filter_adder_mult_9_addition_add_19_U1 ( .A1(
        my_filter_data_sum[14]), .A2(my_filter_adder_mult_9_res_mult[0]), .ZN(
        my_filter_adder_mult_9_addition_add_19_n1) );
  XOR2_X1 my_filter_adder_mult_9_addition_add_19_U2 ( .A(
        my_filter_data_sum[14]), .B(my_filter_adder_mult_9_res_mult[0]), .Z(
        my_filter_data_sum[0]) );
  FA_X1 my_filter_adder_mult_9_addition_add_19_U1_1 ( .A(
        my_filter_adder_mult_9_res_mult[1]), .B(my_filter_data_sum[15]), .CI(
        my_filter_adder_mult_9_addition_add_19_n1), .CO(
        my_filter_adder_mult_9_addition_add_19_carry[2]), .S(
        my_filter_data_sum[1]) );
  FA_X1 my_filter_adder_mult_9_addition_add_19_U1_2 ( .A(
        my_filter_adder_mult_9_res_mult[2]), .B(my_filter_data_sum[16]), .CI(
        my_filter_adder_mult_9_addition_add_19_carry[2]), .CO(
        my_filter_adder_mult_9_addition_add_19_carry[3]), .S(
        my_filter_data_sum[2]) );
  FA_X1 my_filter_adder_mult_9_addition_add_19_U1_3 ( .A(
        my_filter_adder_mult_9_res_mult[3]), .B(my_filter_data_sum[17]), .CI(
        my_filter_adder_mult_9_addition_add_19_carry[3]), .CO(
        my_filter_adder_mult_9_addition_add_19_carry[4]), .S(
        my_filter_data_sum[3]) );
  FA_X1 my_filter_adder_mult_9_addition_add_19_U1_4 ( .A(
        my_filter_adder_mult_9_res_mult[4]), .B(my_filter_data_sum[18]), .CI(
        my_filter_adder_mult_9_addition_add_19_carry[4]), .CO(
        my_filter_adder_mult_9_addition_add_19_carry[5]), .S(
        my_filter_data_sum[4]) );
  FA_X1 my_filter_adder_mult_9_addition_add_19_U1_5 ( .A(
        my_filter_adder_mult_9_res_mult[5]), .B(my_filter_data_sum[19]), .CI(
        my_filter_adder_mult_9_addition_add_19_carry[5]), .CO(
        my_filter_adder_mult_9_addition_add_19_carry[6]), .S(
        my_filter_data_sum[5]) );
  FA_X1 my_filter_adder_mult_9_addition_add_19_U1_6 ( .A(
        my_filter_adder_mult_9_res_mult[6]), .B(my_filter_data_sum[20]), .CI(
        my_filter_adder_mult_9_addition_add_19_carry[6]), .CO(
        my_filter_adder_mult_9_addition_add_19_carry[7]), .S(
        my_filter_data_sum[6]) );
  FA_X1 my_filter_adder_mult_9_addition_add_19_U1_7 ( .A(
        my_filter_adder_mult_9_res_mult[7]), .B(my_filter_data_sum[21]), .CI(
        my_filter_adder_mult_9_addition_add_19_carry[7]), .CO(
        my_filter_adder_mult_9_addition_add_19_carry[8]), .S(
        my_filter_data_sum[7]) );
  FA_X1 my_filter_adder_mult_9_addition_add_19_U1_8 ( .A(
        my_filter_adder_mult_9_res_mult[8]), .B(my_filter_data_sum[22]), .CI(
        my_filter_adder_mult_9_addition_add_19_carry[8]), .CO(
        my_filter_adder_mult_9_addition_add_19_carry[9]), .S(
        my_filter_data_sum[8]) );
  FA_X1 my_filter_adder_mult_9_addition_add_19_U1_9 ( .A(
        my_filter_adder_mult_9_res_mult[9]), .B(my_filter_data_sum[23]), .CI(
        my_filter_adder_mult_9_addition_add_19_carry[9]), .CO(
        my_filter_adder_mult_9_addition_add_19_carry[10]), .S(
        my_filter_data_sum[9]) );
  FA_X1 my_filter_adder_mult_9_addition_add_19_U1_10 ( .A(
        my_filter_adder_mult_9_res_mult[10]), .B(my_filter_data_sum[24]), .CI(
        my_filter_adder_mult_9_addition_add_19_carry[10]), .CO(
        my_filter_adder_mult_9_addition_add_19_carry[11]), .S(
        my_filter_data_sum[10]) );
  FA_X1 my_filter_adder_mult_9_addition_add_19_U1_11 ( .A(
        my_filter_adder_mult_9_res_mult[11]), .B(my_filter_data_sum[25]), .CI(
        my_filter_adder_mult_9_addition_add_19_carry[11]), .CO(
        my_filter_adder_mult_9_addition_add_19_carry[12]), .S(
        my_filter_data_sum[11]) );
  FA_X1 my_filter_adder_mult_9_addition_add_19_U1_12 ( .A(
        my_filter_adder_mult_9_res_mult[12]), .B(my_filter_data_sum[26]), .CI(
        my_filter_adder_mult_9_addition_add_19_carry[12]), .CO(
        my_filter_adder_mult_9_addition_add_19_carry[13]), .S(
        my_filter_data_sum[12]) );
  FA_X1 my_filter_adder_mult_9_addition_add_19_U1_13 ( .A(
        my_filter_adder_mult_9_res_mult[13]), .B(my_filter_data_sum[27]), .CI(
        my_filter_adder_mult_9_addition_add_19_carry[13]), .S(
        my_filter_data_sum[13]) );
endmodule

